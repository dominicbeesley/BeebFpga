--
--Written by GowinSynthesis
--Tool Version "V1.9.11 (64-bit)"
--Sat Mar  1 18:32:38 2025

--Source file index table:
--file0 "\C:/Users/Dominic/Documents/GitHub/BeebFpga_Dom/src/gowin/gowin_tang_primer25k/src/fifo_sc_top/temp/FIFO_SC/fifo_sc_define.v"
--file1 "\C:/Users/Dominic/Documents/GitHub/BeebFpga_Dom/src/gowin/gowin_tang_primer25k/src/fifo_sc_top/temp/FIFO_SC/fifo_sc_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.11_x64/IDE/ipcore/FIFO_SC/data/edc_sc.v"
--file3 "\C:/Gowin/Gowin_V1.9.11_x64/IDE/ipcore/FIFO_SC/data/fifo_sc.v"
--file4 "\C:/Gowin/Gowin_V1.9.11_x64/IDE/ipcore/FIFO_SC/data/fifo_sc_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
NShi6fqnLdc8QeL7YgFKMvdXxJWjffOrerIugI0zz3hkQHK/ClaNYoH1eTp7eu3SBCo5oLiCtAFf
kgeMIbifpksv1v37lPyWEnCHol82Q0ftmFtbu/BH7z+99vXri8D6Wbk2sPKokBAh8/MJ3JfR6tiE
UEoc4dYOOVyn/ZY55qSTG5JBIE6k9CjGoSlSviDni9qhpLIhX8fgPcqSUYHjKDwvf9yuWrPVudJe
JBnKwDWvN9+DyY5KuCb2Wl8pmjevBZKzUShGGolFSucCJMAtE39H+xSDoXFH19qy6RZH74a8QQoZ
shdjWc0/bGpG17oURW1k8vdC8TaHFAuPDSOs3Q==

`protect encoding=(enctype="base64", line_length=76, bytes=247952)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
JpVwk4Jko2UO9I8IMadk+5QCsIiVjlw7DOlhn1cyLz/LfOpSi7BWUm6Pew9kWJp7q60bZ7HuATL+
hClh/lpEY+2Uw1ogW6zvdGHAy6ZT7ojCD+1X6mYun/rRgB1aNGy7uUz6i8VgObPr6mFSc4TL3Bjg
DXsWm/s9XmaJo2zKb1pBI5olK+HoJxuqs5pItlb66fPfFyHZkHuy0qxilT4WjzIKg+roj5NuUjjt
oIBH8AeMBWCynn5+junOMOIP0Wpn9vSkvYjpKw4S5BHb2wOAimWssn9Xt11Bxqx3X+h2c/XoPZ6O
TcFSgYW7pGr3calwC+F2WPy+ys6WEe19XYdO9QTilOSR+8Fo7UxYeX4P1RO4y0e2f0xLyIvibLeU
tsXIEOly5xhxFGrG4B8Za4qXWRqcY6SGt2rYgfXmlvc5qdmqIpsIKkDMSyA4P7HrxJfgf/zmvOC9
nrtnPPcmtP5ispf82UsGfKqTYoWqnzq+D20rjQY4W76IlRojKcJbeWwykweXkpNRGOX27eRk5DQV
bE5kKS5BfkGX5R6UGOnF4eHgsUnCSn4xWerZMBmgnICqTe+ITbfuL8eg0+N4nRzkO1sJxr53UTfC
FoVs1eCB8QYGNZZNOp0NVkREqswrxfNenmUk6s7CoUKCjWN6DCtKjHRz0RF8oJnFYCHJ0BJTFRLL
BiY4xCdq5F2ApSAd8Sx0/QGtQfAYSbZEVGDZOjUIYRt+uz57pIaZyarvbqKlGDeEWdbFBqsoCbrx
sLSzoTHoUiCP/ptc9xVx2HSj7oKv2H9IuPm559DDLy2q2zDOlK3fQEELjKc2TsY235vdU7UIfNi3
D+DHegSgJuVs1Ffl+6ocozl1h03c61l5VBT/k9/KPYFUbRUZom02THo5cpaDF8r8rxgSc8i9lE5S
Gb244iJ5WsQyfPiQJazSoJvIcpijHThPHkHmxUUsVLTjBd6k5zSamC84HCSpbdur2xu58qcuVnc6
DGue83CnPYx2D9enp/XHeX8dzSK8kCOTwl7bvzBZDuwyO384gBB0q4rolpNypXau0LJneB1Ugfpi
+QYS2/lSrZTOclsSdpjJqgAR1KAeDNvrQ+iIjgtoOejvgSIuQ4pG6TscE54gpgmwJUdVHpM6Y4y3
cieEN2VzNluh97b1nNKcmIt+BUeRGKdoy4x8FQ7M2i4xo1RXvjDCkC1zR0dRmoiHbA8kWzNYYgqF
s6vpWXop+zJWaSfKoN3fwGi/UBGSOthF8CVsJVd0q/g0sJSexuxyqH3h/tK669uAyzHmG39zmYZh
4lEiWYO3bbY39swNqeEGG33CdE7qu/9Q2JUkDFio9f8pjm29ej5prGwU3UieRcUeKZdVmvYWxK+N
iWYFWMBsBSc4+0PLyk9vNMFnzAKM/d+fA0XBBVKVly0rLei0KzGpnvaz9uGjWpr3uGx6DYOTHWl+
1ZFcItXBqGgC96MYJ2kBGI4zubzyEw5nWLzcUbLVLNO+2hbLDAzc2XZqBV/cQ+gc9szYKKVXwi+L
ym9RfC5NrPTSWgtS9cGA+eFpWV0ynIhjdCIu8Y2X1dG79NMRkDoeMTDo5TAmwxX1vXt/L8o4hxDf
I2oX76bWuDg++0lUav3PRw7E1I7S2bQPYPVBTkYghP86jtVM05AxFXBVep1VZ/H3QrWMhF49NWh6
Iuo+5pLkFV1QxBEzKRL6SgH7tPVyt+BWz9gilsGMyA6Ihvtdn0VLORqmQzDUhgR9eFG5qgHrrXEi
NXetXBt6G7z3Kpi8ChKhk1pfD+NUQK11yCTSgYLU5nAktguLuYHBVsFtkxZIXKsG67Q762HUMncN
USSX2r5v/9MtTFElzqCPocR4iDXo+61DhZp+s4pSAgANF7FZeuEDoGnj901HZBzYDbN2YSOXS25T
q7ZGwZZLMZ8WZ7FvKw54kQh0VZYogoRWVwcoPKcB4eDuEjm6MdCTvVC/F8PRhIZz4jlg0qmPczku
v1kLt4xxCEr1jWQeUiruI51lIEW+F5iWhPSdorIF0lmojJk9nJsbY76khZUHWfEWu53ncxPtXqB6
3EP/9vVteunH28IVCemXsWfN1hoQl3w95s0+eKzCAj8Mf6i+owGe+SkJxXJWtteXJOXil7VH6zRb
rEmmjAK5B0eGc8/AwRD62gPc2rW6NbhEeAKWVTecv70j8edKWjJG8O9JwYFm/U1wHqqEtX94F+cX
7mGM1qZ+opxfQy5qDLT1erbVt09gna+OgvNLWFdX8nmTXvQOmDWgw5WDlAkF+p5GYB+MGT3BcILy
sD9Bw1xJg2Jv6rDgUEhxAqwHpP7uQJxkQjqSpqlkra4FhD5/KngsE3unj7MaN/MvqTG2h0qPIH7d
gFYAUIs+0XAGvUEny7Di+0xIs5+E/196yKE2qoHHNa3DVFWE8flWMgLy0nmvasdrtEJ2T7iUcBP4
mIt4+tsF61DdQ5QK7bGRdKLjWtM6aGCOI/i179ibihkh7jWAQu8QutZWOuvT1wH6tXfL0NpxtH8i
CcgWVLkgoqnSOhtl6QHhA6yfA4obnS75sBnraBikD+mw6X9lqEQ38XS6r5nbvXZ5bguvPVUJKmoh
gPy2M+hvC7S6+IeSq83M4D2jsCP68kXUjxHl7epdoMdLFA4vmgyypoLw+dIPjdskvip/tqz3y/ZB
LE+R9ifCky/VNALKWHX7t56lIT6uMipOLNgnl+gi3QPLFNTJZ26j7PTO5dUIVhvo2+icq24FBq7b
feYvBHJ1Fyd9XpiTZv4u3Y/BbPmN/IJnkYB+LWXx8s8eO1TRwF5zzlBYnZSGbf6tHF16UIDY53q7
Up3M41SwFBG47+Z2ttueTto5XsJr/ttjQD0cY3FhaLmWbcRJDepvDVUeUttW2KrK7Hky0un0LRgn
T4knaw/8FVY484T+VKtPaW5vkPzGvRSHzIkeFQ7QBgKXGVZvxCnEtLIEVWtcBmubqaqd1SeKGxVv
vEYE3I/Ty5kXyHUVYRkQJNsYH/sGdDSPD4z/Dho6+vLGZauckXUQBnOS73kuXNWip61OeopdJfdC
YQsV9ukUbhff1MHmRTANuH4jeszHLiDttSFANx4M7guOrpA7xAN6/YHim1ElQlsR+i7TOPzbSHkT
VTOqcXvRdrcSkZbIS+Y2nJYENyosBAOr3z/2z+fvUJwku88YNjwDw07w8KUa1aeCpGlavP35M+lh
pyMDTSis025UVN5CE8NYuwr/I0Yq+kyYFj7XVM3ybGqT2dRXX/hmOhvML/qCNbUjnVFsSRRw/diF
ErHX9Kq4l2DiLcPDJiXzbesHY7zVxao433PQ/LmMnduqAOxNljau5LADePiKSfmU0bbxVfZvQjP7
vhtlJ5jZdAI7/lM96iWvZ3x08cXNzo1kCn4k7LHR+1uhN4CkpdQ6+emdccykhnFYuIzP5SkNUFah
ue6CTux5LMCZhqpFkqiK3AggqVAEuI4XyJkkasl/3ljq905VyWbsAmQDYZNxGB2cuCn10m4SwuQk
rO90B8/YvnVJUJLGPRJDnO/F9+OOBsCQzM2yhLeTGbgnCAtDammrcdunlijBF3Xjlk2+jRv8x8lr
Di8w9fFZI5Eyv4oNR2ua6S+e69iW3gBRygZd5+gV+pzDjUbs8b/9ZCSLLKQnChX3dizOr3d+wV7W
eWYrL0QKgxt2XfG1BDr7sg5r9ArFsxjq8r8A4anQ+29y0x9mP62fYhUM4squa7A1G7ooWGXhlzLZ
2hG/fVozkPRXf48tuCXY3RziSRVgL02d3ZoPVSLu5Genzn33n7oR5acvbuAe04Slj3TCyirEa1dG
OoZLBQDIWblfuQuvNbLIKL/w3mqzzokrenxYpA08MPjGLW6IQ8dHT1V7LW/xuO//fls2kaVgiSZS
wJGImal4WPhXcflQ6rrdRu0cnQTkRTNWf/f7+/HkhMTDJwkGZkprHgE4rW3K6GyNiio94ng03FTT
IREgEwJMASxgBWE7dtHkxJZpXN1zQJ53rBB7D5z7bfmwbAID+5sPnYEeLk/Ju8G9r5ZrMDzqRH/Z
JG5oPE6BbO+RzFpDtmRxRQ+puYpdaXVyMgU2p/ugn1HL30UvMM5RklhQQNUhQaWoy97vOznzGBtX
V6TzD4sKAljiIcs9Cx2ExiVbcNLq4UFd1rA0ZKysHhKElK54cCRj7B2pG3sTvvQ8KYUWw0+1rOo5
aRM+IbhjZEOB3LVp/RdPl/CLOKIEN1YJ6PPgs4vdJayec3GqJC1jBL1YInIL0EiRvbM9MOUxIk8X
oiki2++KEnMPt5/v2mYmyFTCc5bus6AEyacMe8qpopdJFyeWn5kLqrWD+qjPHEp3DNTJKEihTX7f
+U2y5Zbxv/Rix3aw1iKQcLrhPSJ8V1VIhCNuRdA2gAnroOrfLOXEcXsZcFMQENf/zfes3ZjCm1DW
mmTUE5oQbzjaD7jDZpyxjnkpqyAEFKffvBjEdEa0iaEYeX9X+E5b6oe0GPf6GY/lscUOhPmg0C/A
wFu3C5wgLV0aZk0zBKJsc3jtums3ipJmFRszbK1eWUICQE3knVjGatko9J9qZV2QJGG5XijX0jxk
y4Cn3kkwjg4X7kNKyFyex2vCbzi25Zjt1H3M/1pA7COn81FgDQbVPKwGiU++gdpk+BU2dLi5LUBz
8JUuIaIBTkhTwFS4+ijyMmnLHv5tJlnW0IYJ90nLr+GN0kIMVoqqCrdoiwJ2SyuaP3RS3soQTuok
pLhLOGoBL0OFonQY4Sm+S/nXxfaLz87CTKdpVn0fj8+KW1r6UpYiT1U1XMqgvDDiPicFpb4UrHpV
pqetVK2lUzfWSM7g7y7uMrfmj8KG79Ll6PaHZOMPJLXQR87zzFJARy5uJrr9SiZJNz9aEyudSylv
8Hh0Ij1kEYsNa+4v+3fQfa/sck6IvdyHkcZco3nIneo2/tNrvpbaYWR48xXO9WtWAMgtt5FpJ0Kc
9uvPPwzpub2MaEVw9Q8fXWLDaOiB0M5/tXeHZRvZLwzrirr/CFrOHmUNGJIQUpzw+w9Co+CpcAeX
jE9Whqihbn9BxMZRAHZdOS/OkI0GYtkiuSWp8rv4ha2da/+K/EyAby0aKK2vh5ZLgSHFJ1PBMdbT
D+5XyxH4PfGdBgkr8s3WOSpld4G6RI5owieZ3vFi4uOEq2rdmJfT5A51R75Ess8GaMWfZ6XrCBew
h44bd1cVvMAo+4+GFPD0pfj/tEfTrRhmST31LpjjFDHdKDbHDZZ9xLGAAupU4Sf5eIlVVC987s5D
kxyrqn3D0dst7FoFtN/uqWpCl+UkSj2xfoIne0rgh2muRHEwX9mihWt/jXkPJoGSqOvbGJo2AUAz
T2e5eIRuCgikEPgdsOpM7c+8/5EpePS0grtA4PGW/kd5nLnKuSOeeygAG6fQbylbY38ni81hSfq+
DdGPD38e6GXImvLv+0davcqf0Vugz4OOmge1DpQ4lJMhk172b2fuqgOi3K0aNrQTgIXHMhPD+y30
l4uhIZNfR5T7q/C7KIUYKly5wj7vuS7/J3EH12xrFyBaDYeVFeg/jTgGZQyo/pCpjspv8aRDL9Xv
vK58SBDMwwT3zEquiM97FqNWvo1nJ1kJDHGjw8ZBpx5uIyv/2gtf1WrzJTmMffqX3faFL9JHZY36
Ugz0S8SJv10K0+xSA+V57cqCGSUePC71juY3t1A0VV5k1Z/1idk/X5lcVloyBo7UlJIy6ekZP1xu
4leUfl/11ZMAKrXHvJm+2f2WBEpkIx6a+S6r7ykden59zkUrcX4Q0hLZLz+8Uvoo3Q0vuYZh1jJb
eekyvArvS9CCSCG+8oYou+qcL9ZaWdInqWFlBitNJnpNJ6RWpCsZGudXImJuvZG8WN5AHfkOBL4r
kGl/oZ9j9jYy8rRZnIBzLs7SUbplXd2cfAkmWThYsAVCoaQliQKumS3HieuemXk/X/phGFR5pWcS
u0C1YMwvSvqIRQWElU9ZDNceLQJCSWpNEGBbgZiZjTD47HGaUXbChioFlTdXcHcvffgZ2lrFAbY8
7F9/N2nsno9OJ2bUWKIkxjsXQsG/fi0HnCX3otJhLtKx8HBKzjY3wADxmGRIzfKr3hkKa1afU4h5
/p2oe/2pg5jIfMmuGodgUwKv69gGel4EpRPIPHP7v8+AqBJe5JSnPU37M1omN+39PupYgBJb5XV2
0HKeBLHSwaWBUX9Eb4mJdcDS0tm90HnnG1Sja346khiPab7ryLYQqqrdXR2VZqbqhviuLmvOB6Ba
KZlv4zmcKKmUtNugdmaD1u5dABxr5RHSX8akY2tJ+L6dIy4Tr7eZ9FcqGDSwiC8R53U49RVmx2+y
nVIIx3LHKLpvMdzvUY11n68VWnS3gEpazGHtN5zbIiNhgwqCFHGHhqNYP9hnvjlAHkKKP+adR6TF
ljodaK1L2cFuzz6Ps4inAym0c90jaqeZVtWT9R4VUk8GA24AQ5rdBtKkRDTMaZOK8DZSokHp7/K8
4cGHP1g8iGppIbO37jnQk2kbWz4ugP5di35EXCkQAT0euETz0ol0uPyXCPYkKnrEJawK/QJMdcYr
cpZh5SssnMoH945dnVMNNdRG7PSZ7e3WTvLyNt1wYrgGsghlM9ERL0ijEI6/CJuizEVUU6PdETDx
bdDNsPzuuc9MF40mO9mLYwLkLAuVbYgUfD7uQVw9jBxzi0cjnj8DzLvp/282fFtR4Z9jmd/FOoJ1
nGLUtZkkj9vKxfgJH4WEBioM7cWgncjO1jny+EDKPWvI/9X0gC009qbqWdbTuQlnWvH2QQT9thxm
WewUA5+reifEakFr8QOHj7BKFkz4yFWfUQ6uBwBrPF03vxfIBNaGkNVutbgbCSABCRhC2L2NEREp
GDy/tP8hgJMFHtgLjdVA4kvT6EU5J7rOIbF+R3XrgZIL1JwwCPnyAG+96gwFV3MZejGFMAQbGqxy
gVa+XwOtI20Akr08i5Vq3rgtFcYbCkBeCAZB2UFfeUSXTmYvHoPbHl+HcBqMIpfy/eeOgGfKVVXq
hWb+/x7r5cm5L+kf0NRbUYBzZSZAx1ywF4PaCasio1Rg5kRoV5BTgjtZf1Vuf1uRX52tar6qUvgk
WAnNzGFGD7AmHfNG339snyHQECq/V5UldomAvQtCGgreaYtme72aXTRZoQ3CY3NU+AW10APcqq4K
Gc7VA537Y6nB+wP3pwng6yADWVbYrs+dfVjNbhvAd88DWX9FsfTnHxxU7Wb7lHcQDi1kwqlDeEaK
iOzlB6pNzQTvSeNxVptLAzs+RRNOstVmgDYRS+ie2vTYm0BbCbtJLr4okPIvPw+ORr9ifz8XF9u0
H9lWBjFj9+wGCTz13YIkjjQkQJVPbdgQUk+rT7rpEomQ5EVjgF6Zofo29HVhhwEZZWKVmTQ0g0nN
kdKXOye7swGl+ykJ2xYO8iEZhTXQ3nQfT6tYbkli3OVenINJ/PyYovSXE67dcSl+fIujX+Cj0Orz
7G8pa5GoswlMpShziybbtoGb9lGQ0xTMZiiyy9Ke+5SGvk4rxUE4GzFis+CvGLo/fLLt9Qp6ZpOM
5NqZdEXY5bLrUobkvMINNzZPCt3SxwyYjD04Ao4yBjiyV5JXkgDw8BWDi6fAh80eWeimC6ZS7YOC
n3QsxjqubKnwUzzIwwmcNeYQzZEAvrRNRAiErTKL5vbr0Pt/VWVC2Kb3f6sDXB/l4M3o0lVlAO5e
2fKZgKqYv7DpDnqxjHl78Kvcy7/LVkv5ZncDo57ZrI0vIMA3mhcH883RS6IPg/hWBKSY4BwlcnYP
FJ51N1mUpqICLT0RY8WXnvjPWem6Fk49e/VjGcry9APME8VU+2Qn+R0FHQbeZLiTNlIidz/ci/Iy
5+tDMqY0kuHrBVBFgI/mmxX3CqiCEpq+6GX4jiyAoUGlK13984aYoKm8aCCiaAOLaK8CjtyClLtm
Uku69ixpG48e/8GZBxZ7t3RowrWRDBReFSx56u5SWOnYDOXCfNFZmAgDcIlX4myDbqdwU9VhLMGc
p7hRoGvGa8xf/V8LZRWVl1YbFxRxegxfi53tmxSiORPVyCR7+yxUHpnDkPQLK2EiIm+f3eEAmLTi
70cYXo/BQMfHiFXYnPrX4lvtskC6DeT9zHCgpdXc2zePmGY6hYwij2PnQQNiGXlaN5I3L6CIbpcY
8791DcTHqtDR1GL79BEbK6logLPPHSv8ns5DFvLTFS4r8LxeWKq0GoQ20I+Kme3JdWcDrYU4juh3
E/Rn0Kjmp0Rv24siwS8h3F02P+5d8Dx2/pO0dDOCV2Ct5zHWnu8YSUs7OfHCj61gprghC2Mx+aFY
AvXgropFyH3V7pneGtaQD2iYTZu2HkKPwDW+YHLGIyHKNtkDfQVSVe9MtXwGTXYzKUON+0qRvol5
4Kmt645ajjhzUOZ9Yn6aE0fJ0JDnHQgejAzibZk67Ps5/DQosojdBMGcRz50tkHLDujG9Y2p/lkR
Qpe+aNNFLqfZ5oQPjqljrqvDqL3jsHSg46MOGNzHtzVyiuJ+EwwcMjl3aZRuQGCOqEWu6QMmqtJZ
5kUwUR42hKnmVkbCwheGKGDz0OJ1wIaaqX/ehShFzgXJQhCe0MBKJUXg7284pT1T5P1b5bJcqKCR
/+azCcmH9psQrQ99N331eyoZyZX/e5NVoAkSVjhMQgt2EwsY0xbEHdCNgsUaL8JKsATR3pxbNwr3
xbEMvT4RKTpTBbH9qvEWp7stYewD6T8HdyGVrkemLu485yO5wE+Iu5I6hIIsRQGgGI1WF49DmKcl
AxZLa3IyZubhSwR3+d6mIUfVq/DODir9cj4btTxv1s9O15DuD+xqGE0sLZDo3uBeMp6hXWcX5Fg9
qZi/CrXvYctjfnxskx8QjKYdT/mwygtuSMfUv6JU1Ih0D7VkEC3GShaZL0hOxGiFy03r973XPRF4
LiSCWseWQZG0INvVPZXyNx/mz6P5TYbEksUxEASzqHldX76FLXWstABOgLMsdg03xaceAG5mU2ei
fbOVP1XPDZHCcLN3h+2MMjgoXL+hwTJP18sQwlygiIZ6Lx3m9oWte73oSvRavEcphtsHbmh373xy
bOJ6uoirxCUpC7phoHBkn0yUGDb+aEg3VZALGdQMCL9EbVhp+HG4KcI/x8+vR1sz2ydgAtIWOd+U
Zw/VasxlOaMKMzkpIZIflGLLfhbuiW0Rvf/w9OUU8oeswMmfB10QpXR1j359+kKsahUvB6+s5peE
2fbcWqOnlDp3m3QPdZtx2VsB7i6lLjBSdzBQLxhNLiWbuyFAbaC3JVXL6X9yNE7vsllv48TKZz+W
EqSABSn8Zvl1b4SPjfGfIYc1zwmoj2t+4reJH9XiQVs9Jh4jjkkR8tAbwJ7r9cRDEsoAWj8YdcEZ
Dr3mF2Ro21i+OjgG/a/6QuDJbVVqQnspiCBoXBSb3f4pPDmDKweo/w5L94mrE/VzcouvmL8eWM/J
uHLThIdTIkUfFiv3BHk44Wlbhr0tXryNatd6LQFiGIHFPhFCjCEHaeMlKMzd++bRl3NoxndpMPjC
CY4aIXP/DVGbyia47d0oxdCPF8uoVH0yYA+bESICw2l/loWMgKP8DEFEXGo/7WbQdzm0aCvbxS1a
jD5tzpslXw6YUqFgNtAwPW8PFvA6jxpMhGY5Y1x20nTdRgg+9fK8ySFxa700fQLONOzeEWxJlZ6F
nrthl3Xs2JCVasrsNMYAXEpkcUmpdL3Ai/zrzH7RsQnv3KC68B97akGaixB7CVRTWHdQPa35mpoN
5tqHNUNEWEJhYB1MfFROyt9OCaWitDmebUaIju3z/rzChVgX04ZBUx6FjM3TL/mGSHZthTwQyCNh
d3+8xVqCaxWBse4Krt3Z8x3sKNx1xMO1Rryy2c7VQWIeBvp/J04z+uaPNyiJcvwCWsLIBU4kJ8KA
AlfJ+Ta776EwkJ1B3sBKaU6d7uNPU02CUIK9xiSr3vuNXpXGPBsm3dj6AAbEXBYqFfHSqawN3b6F
mZF42UGbRAcsq+DNOKjXww0CxqyFrLkBIcrE61X5MhcSjurK63VoPhQmG9/+aCtcnBxbBnThOYxV
HZmFVT38TFFEp1gTfIdhke21ZpZeFr0STH4m5fvbDBE5abLRv2DjDdySY9FK3nYHutU3H1i0HryU
g9DUABN1uQN2JQVq5jPRkMpgnCWRffuZBBmkWoX+6gvV75HWqjI+fsZIfVGvvTODGl3hcZPxHnWo
GXhxcxj21ITNExVtbVjw2uChcFVAddo9ThVGPyZkf4FFaWunN5gtqTp//1wJ8FKdNMSy4+1PMwh2
ymfPtiPN9guvjMVD9fLdtUDEAt5eGmJpGxI8DPHMdC6sCwOV4XAclrQi73CZpc6P40S4E4XRWJOY
74/Ow6tmOe6aG8BHjGYWEFcgDetIEld9nBcrlgcno6/2H/nkBTRdTQ9FGhoJK9/eGkKNs2Q5CjRX
MavxKpxK/JldF91aJbl8uURr/zpO5beM3ZMjuxkNGJ4F6yFgVW2j2GZ0kyuXORFINt1LwyHPJ7sf
mvrtFDNC954pNBfPn0A3kj3K7r8E0cl61WXdsVXK/oPUDkheWHDbfR+THbdYUTx0Ib2Y0WXl1isa
YV0ZEZp5cvibMsV+adDXggRrThVqC6XXHTJ/d3+GaIJzHwIeIU+ENfSe6OAuGj2B1/PgLBZTOTx6
EsMhXpERAnHFJqzmV5zSYgF43jpj9MveS/z3Ujt5axtLhtumX8Ta9xXyfZdKKSgn8liu8h8e3f44
rGEIv8wlZLWlyROdUyXw04rw9mb0tL3BYKDL+zHsFeWOT9LFVwFCMQyfqrLU13PxSSb7nau4ES7U
xEvZn5b8XpmwvcBbq5SGnSWPLeWKGUGK0xkpNYSL3bW0I63WCOzaGoRwRd3ANKGHRnekE+9bjsXD
hYTyO4PPlrioF6obmbm3vQFjjodYcBJ2fDW+LAW5gKUPFh+TYgLyIhEXLz8vkl/yeN7AaDMClPSE
PkHNNAoSEP2nrac60EMH3mltHp4nQ1cN2J2GhtrCQXIx41c8qf/JE7WntWAGNn7eE7wOO+JHxoBZ
5tbwFdt0QVnuymqcWD+cEAo0A9mDNlC1g41nI5F1j1yQuFGWVggfo/klBwxuSztwUWXgUjB5tdDL
5+lHUDU4GSfnuWi4k0vqFqP7+3n3YREffj6N4cVsvH1E15n9SD5qkgQuRpLD3Yu3PZWCVjPRJLj7
2i6EUmpoaU3p/TTkNemr30kwILPQb7XmGYcHLMH9WgGFzhDpMnao2wpHcuCw/0A81qAYqOcXxBsC
L7MLXZ//fqVkl5YljiNDl0IhD1JFVzlEFGOjXbiF/m2MwLbhNkQ9BMbUgxwEG0tVggN3oeerkP1A
h1TFtE1DEiDWvgTJFpg0HLXIDBw5tbGwsm3Z8G53bIjiJotbr7aapujYzvo6H9jIb295LCL+4FRB
vxb5OpIeSLewz3hlUGpmV9TpvaJlDiP57BbBX53TH/JLVhn9ldEL8crTCop7PEd17LKNEcvL9kpc
QNLRCjllQSjVjNuIvDI8YsfXlkhM5Cwg0DYnOTgUROtOeE/PBOt0fSOwDKfoRvrQdgIDvY8tHGVf
mWD/0B4PDsmJMBXTi/CiAbwx2f0jgAxIzt2xfDacwvkA4/Qg3Jv6TgIneFiEJuUWFg8B3K1ZFIwP
gu5lajez8i7PfOyuvlilisrUAu8lp+pbN/NHAlVS6CDLmilP3MORJgdw54K5KewKpOo+0d6SmOB1
jSP5vMwagg8vgKCIab+CjS3Om+cUFUbxpZJHJgBqEM/V0hCKwHu4gDDHuwjIiOvmXOydFxwT21Tt
HzZLhh3Tvl9n2Wm/4CcuEsxEBRZS8VsHyQZrLZ0DGljEfLs2LKxsUrAOwA2YBzTaXiGYC5HLjGV0
JgDnztSjPx5fOAfWtUPfqyIyJs1Tg0TldwMYick7K1MknH+bC7nb88Kn5c4P3b0wXH+nBVGVPBf/
rz3uC1NjyGqAJ8RaDd9Qd1qbBaahdKXkiZPt2gayu/6hleM2yoRg6jDevd+/MQud8uxqG2et6/o4
mTAfPtNrgpL77UmHqL2rXAtfop3VG9oJZ1eXcg9m6bugK5UOrHvap0a6JUE4dykmHHiuQL2pF+sA
MkDpHZynTY/J48i1fxCV8P5TNa4OUtTXU8QxUuCJC25N+DTfwyq35ifdh/yCYQpDV4RWUtQJHJcZ
cOa3MBbJDV85jrU/VhXZzL6k+qMKK8vZUTZs2xpgIFtJyOpWJuulmDZbydkp9Iq7cNg9qLmc6IDu
i9inPqW+xy5pX8skjjySqXS6SR3Jt4idjQcI5JTS4NCidIPc97fwlsHwqM3jonuP3+nIx7n53T+Z
1Cgq82yavnl7Dxn3zqnJiNQV/5EM1nyuwiNd6/xm3MwuhwCwycbH1UX/DFgkrak/ECWcxTzvAwrA
t35PwVLznh7K+iDNhjwH4frBQctRtpp3LultX9WdOacewA56Ova1OWJhEhSh1RAEP202QcZXFee3
D7UV2aGgrt9v7Rwrw/+ys+NSA9U93jwAOc3x/qQQwANnG1zSAMfaYsoPWCA/KefIdSpcai8oz/F2
E8SpSKS3VKo+63V7fYSv9eeA5mZ2p8qgj9QNTheLmaxedPxM2lnHZjizBCXQ/SmeVzIB3vOtY5Lh
iUNuK2gBm1Z3VoNQA88zusZger/O6OaOXBHOjoKpSPusuMvy1qQ7SykvyeF4tlCt0m2h/i8e0dEH
Bks1lMUwirrDauLoawuxiWs8ZL8C7QItxJZ5j77JL2x725ttuocdOhD7wnx7nAFjFAtEKApXHbUL
MEN30KbkuVMzu4AgOXi/S5yH/M+y/KKndMCk6GGrnGi1/0HqCnxpJFqxf660N93uBcKadumP474P
dYsmDUXGgDp8juSNUmOEoEhW6xk0nlza/gXBE0GhCckdwO4CWdC93q1V3MrVclb+2mZnbJhkHxNI
ih3oQzSKOQSRpT064ZVHKsoylRKMecxoI2AOl5tFDBRP0GUiO9T8X2HLX7tqcC+NQ4nl+yO4Qlpm
gsGkfI/aJNqL0QxVTcC/cmFqomzjNB1B8knmNH+wA0KbIcKpglkN9n2nAvHRfPgC7Opgf2B7raXW
GyhcJxS7t/FO12/5h2Yg5lot+8n4XrM2ejPuHHRJccdcCAKUrkNfRuabnIHHbDEVStuiYt8E1HAZ
ScJ+ulXdxc0PJkBUEQGBIfo8s1SgF9x0a5FCAUDl5m2rYgT5QuAMu0xA1ims77Mwf3hJzOr0gxex
+kXZxT7L9yajDsKG6N5zGsiUT3IiolM7FDEmMkghE9+2mZXsMtNeMSSkDR4ScDZhX3ftV1ovuu5L
wUyaVs3yqVuw2CizCL2iwyGjmhvAxve7Zyewj/2F/KZOhy/n+x/T2i9k9HL6HVx/hp/s47y1waij
2nDosceaD8uJ3qRX1JWIMEFEIQNtgWsL7XCeP3Epz5EIqAQSaciY2jMxDPUn/5pKhtAc15ufKDml
pR87S7ONQEkjhMP+Tjzwe8K82PQ6i/m2Iem4FK1uXOCIkbtkJECe3Y0ZzxH1gd2onB/Q+vAH2O6Y
uAW3i7/w++xn1OkW5OsXrf4Nk7nq7EiUIMNS4hr4G8nD2+WNyh2l6W/YMKzGG6twgwtU5zOQ+AnQ
9IoDhO9X+tAx/lCS5u9IGFOLZ0qdqdO1rmcEK6rMO/Nh2NyKo2kHg0Mn6zRglsZKr6KIQTiY+AXi
GPcjtfNowExtM3WXu14Q2KSi4c1A/QEiHl6lEnoN/+wmFNA7Oz1vbTr50cYM3sX8NOq1fTSHSKi7
wZmrIvpYfIXsxuS8Pv5wFvaoPQ73phOQg6htSj+BazxQOdGPx2k886FXftBIUELJFqcewC7xBn/g
aTsOVqqB354BgPw/0bmKc3FPpHJONycpxfSDQ/CXMPiPkild/jSINMOlzx0R9B3c1/faAo6e4UAi
1B35H9kl/J/M7zurjB/EauF93JZOk0YRMg09jSfzDDavYiT/KWF+DKWs2yBCVb1bTz4XOHh18+Jg
3ddM0vQviuMC+1w2AWC838ubF8aC1TuTp6Dhj7AhIalglPZ0QtCRxV/q8/nf1PtcIMEngv39KNgl
gzSZs3/OfjH7dN/hl0wFg+DIx/n0xFmMnIUynfZJjgr77Nur3I/Yb8YyjpBdp2qSW/XARhfXVpzV
xTsS/o5TLOd7qT/SVR4kqo9bHH/iwc5XJJWG98mHtNT1UO2ikET6yAn3tRKiRGwNjxQVW3MvyhL8
sGpfOXs+lgCVHRGbNhDwEdnq4XQ3T7JFNkfgQ6Jo08KpTiR45oKB34+q8uCyG4ffeIKnQHKNyfhD
NrybHzRd3mtHl+Oun/LJ2C3fC1OS0BqSO668d3YYYqWYS7jMcwQapeLSD6uJjgk5qNZj5zdrdJPv
cTbbCLDFE+qnjaeaclMeCLxbUoySuWj5YicFYpn0MwUJLDjY5XVhjV1l7FTjYJVWFsmtR3KwDDd5
HrWJLKJpdP33fMyevd7nusyOzpXKkFLTD2+Piig3dX35uMdVT1sCR8cWrAFnx6+8tNxte4vxbapm
CJyGzNAhNOmlHinzJK46LGskC7COnVScOlLlhWKeEBEkTUyLAfEuQJolNb8x5MG6ImYuCrWkAiC/
ZB/igxKR2RJBALPQvJoUXkbX3AfYJHVPdAEwXGTQjN0xMzw5a7my+olmhqlI1zeCMuUaNpT5U52C
VzIzyYR4iCxeEPQHvH2AZQySUDMSTEG6eu1G+K1C2An2ZdtbHSAUm2vqavaL6stqZH0wvVUu6xTc
vPB9VQuHz8yUqaxruV4uc/2sUcATGze9qO8Ufihv84r2ff4ThNxU7M73C9snS7Vljz9ymmOcVmyp
dhrtmW3wSUu+utuYTTHkHSGTGfaDl5MP66nl/NvQF3dbozPqYyQSp6/DOAnzuf98HglUZW5tfPqc
ns0d8FyRdG81UJIwJxWC53hz/x7MG6Cxf52ep6ogz3/PB0ULQveqNYBl38iiVU2bGbV2UL1Wbn24
/zooGPssTJ2DdzVb5lWhZf+U/Ny0xS/iNeJ4kV+zb693coHObe979QKlCDC6OzhlPVQ0y3yMevsz
rzgXbduhEIwATWBnAbDsOr8tCQjPZMWhvYqUkCSiKYzyRdeuRf+HXOVK3UcgXZK/g1vycZzIvUUW
aB75ROi52aQQWKPwNjoMMmwfVOXcP5fY2Qav8lZMnSF5e/w3GVQUPy/RnjmQFxO5vSt5iL8yros4
pCjPhRIcW45UmdyuWpuyugm3lcQDYsYpAbHt4iDQDoKsTa1+yTytUCfJMU+Sd4JlGMXgsYNS6HdA
TgtK41jvFgDKX/sfSorvjBylBkzBadxyyAjxEYUjTU9dl2kIrNQ3WQ6362UZPiryyQYDvRygD9z4
pWC8wgYap+sPI3Xw0b13Vp+3qsu8rcdeId5u24ym12N+LQ8N7LcydLizAOnuIqiVovQ5NZaZ+qhL
MAu6oqlJztZow40zJs3EfPCXWuIhBnqRC3jy797tV/ewvSUi5Kw/vEH4jNbBKt3y08SID/6PoxPx
gCoAhr1YVquS7+ISJG4LUIJNcqoi6kDSPwKm1sUfTRrENwSSXjhZwdRk1G3PISmTnHUh+OttkylR
2VG2PAW2ITmVTvIsyHejvLJJBI+cr3Vr+Ra+a2L+rflhUyslIVtPiTBcw4oj3XKJWq7Wl39hYgYn
chl0jL4rkB8WG1248e8O5WblWsVoZk9Gap7mqNb2g1Ce/OP0++nGthFM2nZA4JX6R/wYZluD2e81
6YIWm8ywNdjRDnWTApqhdxjjfzbLM3DWZydoJEhsG3+N1PnyILdnvP7G1WaimzV5FVBWkGhoiSTN
h2Uz/XSDEXIpUEEIR3v7qO1MxjEDgmM84YY80P10AJ4+le1MjMOix1XESkJN1U7ksgU71SblHmU5
Imz6Z4rGwmHE3Cy09S+v5SeQcj7/LAS7Ez+86psE0bNfAD21kSW7SvICaXx7pwtan0olfGV4y1Zk
DMHefblFDtSgzRuMK1DScxZLYuXcZihzwUGTXe3Dw0d7YCsbaaozorVfacf7wd0UIxt15wZErAYq
Bp9ea4eFvf7LbCUU2YvKwBCiokLV6iPXVdRR/tIOVKEgHBQjFReFrDV17bcw6KKjDFzF5jzawwi7
DiaoUqUyz1Am6nkv7+H3q/htUV8LV04tvTJLPkfeW5DDZFpyW58UNrywGf6iMJpR9t6jQ96VJVon
jLS7n97xsdDW1hgQ4I49SMevWTgCNbTd8PjO4YgBxVtcu693/Jagf94bkQFGyUdQzw02cddH0S9A
9Jj9KAVXKJVGSN7oy+dRYoSKh3WCLJN69qk6uZ/6TC64dDXfOWpYUTaYg7TogbhMBOJoTSIJjAFN
3QSoHND0gjZ3qjgugW6SrwU8Jn3LK62o1zo6jTKf8UgR7QcvjlnRTV+dJbsdm1XL6uWW+XTCJeq+
3zob58CMjnmK8bFbOnZNe93Bd4J8WI/5s7WSH8Uf6UnMOpkVMYJw8KJm76WoSZQjHD96GfHp96ss
XBxrPGxbD6HWfjIaA9eJWt4LkIQo9kj2VImeT9p6qWYPoTQIzt1i92V/2PjweALvUDDRYm9UHRIy
SbUxakSSLHPm7rWW92Gz7fMWZfVhbfL+u5tSPWMPh8wHFX+u4/ItWUfUPRQPeoScILf+7LM+lI6O
IIYZ7Mlihwljai63m/HCjwz3Su+JkmJMwFdPmS/TKXyK1/yWYEQTols+Y1peUOycRUTXjrXvV5NL
CLMzNf3se7O1GbUzHqu6NTIKOHWvJBcEdhQwIAa3M1IcwbBCxVf9ijKLVcpu3ISmYO/Lv/VR1MP2
X80IoDQm8kNkO8oBlifICOSGm9Tab+8Dw+FK+j9A5Hai0/0G4797UPSVxgbx+PsqdxfE9wLO5IQJ
duMXJZxCkNOV3XQn9S4MUbV0JBnT/aQ/15ONQ1cQ00fA7JbsNtRWDBZyuLtU5Xt6Hi2j62iuFYqE
gcyJFQXWeE/tpDcdZt//iKwZJSTuR3cw/Gmkk4k4XNBLmCD0cA+Bx0G5IBusrNqpkOx0MfyuTMHp
oqunyeiltaVbVdfuEoPm7gGDFh/cACuBo0pp2Tk02cwKrDfN9W96X6HssxpLwkTrqVjz2F3NUB0h
qGlijnJ9KX+/jRogbrtyBW3e0JIDMawsqRLvbDFF7CY8mFroHfOerRf9rCXUgUYiRm9PSFVitcK1
+U4g7RE01EXxrBXhSQ37PoAgj6uIIU4f0TUJ+PCUaFHF1Z1Wo1sqA5eS6tKSHaTPQV/hwIXVGJd/
4qEARyIoi4HS8mxTb5RL5cEGiimrt9J/waxGfVdvwRnLCimgXvlNY6iOn+jH+R83QiHslsMw8DWN
K6NyBnjNSdP3WGStoJYQQ0rxkIqgYbH3ny1kInk/atuDQ+7J9we7Y8/o8hF6VIxtfTVy/6CjCbCw
oW3aMpKfGISgXH8IolkbV5jClj1G2ae+2b4ciihKDEeft3AFmUd9sbBfLOA0qwRpoBcn6t5gOb82
q4kvo/COrfRvexrvLhc0rQ0QISyzg48+91YJJrODDKqw4I5azR0+ThLgBLYRz6BVbCSSWm8Cb6nT
sJZe6zK/kDKvHS07WLyIFDtP8dNIxv7KolfHfR/TMncHxpN+6Rl9zhpcswsPniF1+I4vhK23NYJ8
YbQWzA1N98W/Oo5WRLuXlyLSvN2IPzUf65dzgdrL28nyG7lRMakWOa+7Jt1/l29HFoUIB3O0KKKU
2kf/ly+7tSnOd6MYz5HKe+Inp7OrnC1fd7hzkb4RrMBmZkGo0R9WCKyfx80s6Y24YopsmxBPsnSG
Xp6/8MeCOiV140LMH8+Dt6nelZRimIDK+ohB7+pjkGrm2Ov31MW/GtzQnLZXhtVY0HRCbXRijHhT
o1amL7zqc30cFvRWM7yo6zBRkcepzdUqlCjHhFa/wubeOL7Y9+I3QmoLbV3/8ZOozZiuhVN7qfcy
TmOKxU3/Zol3L9GPrmwI4HeTS3psZmFzjju+injY89J1mV+UGzYHU4Ufway9SCWVl5GUIw3+a6hJ
z2MueU2oeqEDFluqIjO0sjRZlAC42vHTig8An5LX/YqlMVMV9Yu3xK+S4hfPO9mw0eYd/23IvAO9
a/lIFgtCizUEIegEXswNta2GgSIuF+h6H0xNvVhwH/2hxIkt7CqljEImNUUY4bHZfaidzDXVd3QG
fzZhFeA5X+82YlqthO7JYPYsMRE2+y+5NsiueF57bl64ORe9dTBTJ4kzqgE9ficIKVaOC+gaR6/A
BkNDw+oSxgmaAIiRtW+e2AYSMGllO6UNNkUdCTWGH7cEg/V+huDkiYC3IBwgSm2Ul1RMB96QFy1z
Z/qzekcqc+X7bXtQVnKCT6oNO6cq+g3QBW2J/atZoRpfB+N7xJ6YREhWiU2t3AGqSDCrTFmDvOuI
vH7ZP/DZFSvfTwdC4nusGPt8ioeipluYKQC6vpAOjZDe7xwAfw3h+4Rf4o3xa60jK5aptvQQU3nF
rLUrUScobsq77Asrne5ngQLN+CTEnGx/HbSAQNC5n2X4JgaCItUhbJon/vpFuvypD9U7cYK5WSIe
xecTYvFn9lMThRcPHphVVbyvbc+mKCnY8BccZgA4yPz9foOTOa7LXKR4M8sZQwh2PKwSy+HNdBoG
uFIWs6tnbSURMc4uITM3ytS/AYI/4OuGpqXSSiyiR+02SMbcCSgEcpmus48QoPwAQmoiVaRk9a0k
/61eZNr0JTQf0Grjsu6zReF3/dCAluS9QOoA7+crs7hDx1ocCbDnYqNkvCOUcnvTcrBBDN/no0RQ
mFCucltIOatOPkz4mwUQYvd41c/Ev4P9auoXzkO4/VwfSDrQqBbgDEcfPOvI+5KqNR4ZQsnzvozL
F+3rhCiPU2wU7/MLndROtVzX8ayKVwNDdq/4Ufu2BoPeDl6YwEORmfkNubxTn1j2gGV/yi3SoCHb
SWUo7pyRNk6VS0+T7bZ64CmbJ2Fko9m46gEqFsW/iUoHbJDEiFR9EzqHWM5lMZX/lvT5C36CaaOc
H4+BbwmwR8mDnfcq8J5l6wH8M1/IrgMApYIiLDqeXtc3F3+pCgCea/wD8mioq+fiWw+FtR9vPkxA
yRuacDPN0SVUr+q6FIYiTFlAVayDYZUcwYZ71RCZcDehXXKBiq/C1O8cC6ybttsbLlNbGy0/k1cj
cJNd61R/tbbC6AztpFuwnbDiAV2uOLdGAk6iXqj4aaqy0VKopRI2QawT+Bm7HGl0hMzyB5P24ePi
4ApH4wz917Socx7h+qLkPelRslg3NyFDRvKa+2Kk/fFr6I4nfhEiLNG869wqzT3TAAqIymLX+nQF
mEZBCitvgbdebBWRkIScTQBj0Ee37ldEJUZT2Z23k9u1F2zUI18Qr+VtIC3wJcDdPzHm3pDIy/Hb
WsWzrK210aaZbOkJSVtWaT8mtA/kObsvb9iIS7p7vaLz8VPWAHV/CzsGCS2i1grLgwHfsxLV30XU
7h4Mkm+x1WB/eEcXMPEAqgw7puwU/qxYA2gzgXFZQTfHGukOuqsQWEbfpPOqG4WLwfYh6dr4X5PR
I0Dm/9zoDbyaPVF5xWjsc3hbqdd7JhEfhFLu5GFy3oxsFTowky9NujBT4XcG/kHmo3+i6OFOIN80
OitYTGN0bBJMbTnAbYtjJeeer8UbToLt10AYXxVDyolSUJU8pN1Ywmjz1zO7RsVXX4JB3NVFuaLS
kaO4mtBq/adiMSUBDuD7abfJVAKC5fs3/N9mHVFS9PNvIGMxwGQjknQwdA7Gp6uiad9HEIEYJu8K
2nlVAjHeM2TPwKJyJvbMn79+cSXFHfTZ9tvIe69w0xnl0RlFNd7naauBBL1oVk9c4fy9rZdb/lmU
bpU+YlNts5NcddyX3oWO9NZYq0a22tgYuVDCNU+cWsM0rtP0ogvYA/4230eBBCBv+YLANLWhwJm/
HYa3bt0JjJUnaAbeyDQgqQSmWnVFyWCXlYcw0wVW5BX3Dk7AD99nMzzorNv5E5J2Jk/cN6nmAEvX
iXw4D/7bK8fs+DzKGTbTzhNA8hDTwfQ+s2jGonIfRlHIozuDQohcZdaz+r1hBtEaB8yKInSZzRjJ
nCrYSTG3q3LTu4W9LVVN6Dm6m4dE24eghqy8ZvG0aGbOmQZ4Bh+vHqSWLy+Y2MKg9FjfPjm/YhrX
8SADQPiZfzc0axhH+GxE71ngZPs5RC5Doq2+jG/bP662QXsE6FfsCOYENvPSpDKvKBn3UUIfLlPM
aL906BvdTaOTiQXO1K2gEthe/qzTKqbn8/tLUV9ScRviz4N+Ybjp+dmFWEKN4/1EqqggJ+9yEAqA
hUYpwlYhZHNkWoB4T9dTHFCGiorj+vKMHUGp6llrAz2t8RFt7iHTvlV7DSNF7dhU9xEPjA2mo8s/
PlttIrv39s9Y7/9Ujqykk4a/667bPuxMayyv44/jd8i6X0URqzZ8cFzorANjgwQkMfzjeEeyB45o
JBW6KGaVyLGHztWqiUxnIf42tE0wYjdjpWrdMS2RIs1pt5R7HMNySoTLn66DwnQqo6hXein1WACJ
JnTOmfFR9WsITCpX22IlrB9jqqGlwH/L+qO3f6nBEEsBk/aLBH1MWeDXHiO66FfU9ae6ezGnnHI2
NG3dltum1AaRYcdogCUVpubxISGYwQY4UiQ5EhxgMEdnSLBOJEhlpWLmCyab4x+Nq/e9ewKWTns9
lBRfg0ZXX6IbV7++5ZglIGeljBWto4p5mYvS0hoD9AKhZs7XXZYDXuDVDnWNYrqU9gioWn6ns+Fe
bRDS9gx5ZOUDeya/hLYgsjIS8k9/bkiqybTKu9w2ruPlLeZjzOLvwCUZ27kZP5t+3N9NQeYuEu0I
015TjAGxqnbqkZQ+6lXNDeLaLvXlfGvjUwc6Cql+uaoco+zS0Op3yoinFBYtOi9XmJHVPrQ/taBx
BH+B2PnxvzDYjz8ESWAi35xm9SbG4V2cE4d1xpQMkLhMZ3HMb+UoesLmoxrjKzfQxswF//AvXKZM
2DWz6q/PU141Q1wdpp1S+sDGD1isw+MUl1DsJn++0uljjX6U2V5IYlUZoWZ1+PEbjTE0mcdWfVYj
K1g3oz7fEVzmEgpQ55lXWAL3yri3JynJ0TbkGtsllXznFEZ97zMEUB++HYTv5uY5L2T+J9ROORMN
1lq7pL17l1c9HYv6nUS9NdNPawESR9mwloRFRpMqx+ORKqDV2F9wOVTlLxTZqRecZPX3ssGyuOdG
voDtdF1DaT/FlVGDNQsue1+O5BTHCSeddZdyRrysBNKJR+AtYdnlUg/RH3eCavcW9jqbrWh+zjN5
Dlbp7afPheJ/cbSD9RbUKsyQrJ3BSoMYV8z9EgVTYuUoCzmu/5m+0MKQgl8qOg+3dZ0r9bTxe9GW
sRogJwezQxCIsTm+aCan7dLMutOMM51cta4tuoYfWOUJYOcPCr11Wxi7DxI81VOF0+9WpozSPp/O
kCUH4Qp3tBWFnLRonhpafR62k1JMJiXlyTKHk9Plx+RofjYlRPzvYeXGW0Ss1kJTrXTCIBAwaG8/
HME2L1QUS90x3t5V0R5/te28W3CBZxk4UBvWnHbCIcMS6hwIkq3Z0+QnMxJ4UhueI7XNprwfnHtE
WtEPr1ChYafT8URWSO6KPIiVQ2snFebQS4q7DPN35e3llwUSMPRfsDXdmqWgVjaehNXaLS2KuhHm
4uFZnTQUYaF5uMtSYmu5GY+fakj76UKZAtSchrq/qz0sJ0aljRg4z2ev8TweCg62GNCDucgLNrOv
C2Rxrpzkdkl2SwhSBvGhBH1e3jz/q0Jh6OP+BYMnexCSJtRtbS11NEyOx7WldwVyvjK4xpe1kVb3
ZLGjeevSuidhMLnKtwKYiykPuxH2+M4LbXUxc6OoRSKgGPRMKSWUAmin4nBrTy4Uh7WJYpytXjEN
nhvS1YV44/s3rJPaRpk7o2ZzeUbpFrxlnOO5B/pokbVHZHE8A4AJM/iC1Rco084QqE7iwBhUjz98
ridOKlv3Zxqv6okBVNdqKGBwvOb784ehuDmLDU3+XSi7ApTgiOcohfGh+Rs5uExav7/mytu6/Yqp
fvnEvJqpxaRPrdu57gIu/HZ7Mr3Yv7iGhdmHw0S8uO6dFVM8tKtl6LIPAeobWqwj2iwFuSx3GE/4
e7ov7MkW2ujdoC4R63+GruFG3rbd3gTseMOh/u8fnrDpzXrN2jIfRIrI35g2wuGgIvdetglMm6Y9
6f+FAUSH7zGPd1qoJxqZppNGW0yQnpyXboJATJ3c7yD7UzM8vE8AcD7X5dg+s9gCHPDZuIhHEpEO
lOc9KMGq4tRGhkVao8tgvoX919vp+Ur6SLiZ5sWyAf09BgvoznVzc35YaVv4lKr5LFDkY2Uv8Lss
nGvqL+WliWJsAvabd8lAKwGFJShx88WrWGzYJ+C9i4ipBJsXqgd+r+97co08sXA/XKPfFdEqF2rG
v/c9+cMBPxpTW6Cu59jMcuwJ9oSTQqAkV06fCl0TQhqL1pr4MKfI2SREkT6M7PZdC0nbAeB4G59H
XrN4uNMMJc3sGGm1uulw/AvKkuqYzcilsenoH5dBZ7j0mW410nxuq/KZUKZaS1w2/IIArFHADak1
cDvoRA8Np331Yz60jQ9zPQnBajG1FCxSHl416WgZTPyhJr/N8RkIDi0JhkKTJuj94y+W8awhJFe5
Lupp78oK1OGi6zMjdvMzvnyyjlZNh0LZraxX9nsMP1oD8sqRK+6/OGBsnqLHkWr0l/q3uXuYAA/6
GnoOowX2GZpzjDd66HbenPfx389W+KJ+bi6TQ7P4ZOiVmPuSyazBB6awgLCPufdDAau3oR+ZGlBf
+V32xF2bH/dJAi3KfYVKEk7CUCm9mEgVHsSXYYQ6S7ChApp1hfLszCsXJ9jnxRjytajM7F2b9HiY
ti5AbW0rmV7lWdXUBf5OlRboTql2zXtNlPDVeDpVtgT/pHkaSBjHyoJkVwgRsqUNhlHdWgkHnSdJ
dOv/QCWNpKu+g9wlpggR76IR4OhY0N7wo4AzKZ9DcWSt4rqveTvzZQa/3TlfiA4cSksDdWC0DsF8
H7R2qSNO7FOiWiZAtfqZtu/IOwMbkDN5WoGlFWCDmIBMEy5foqk70MB3TmDcYQLfR9tgya3xnkAY
XIC7ab4XVBqL6kG87P59u9JxDoudF5UvZ52mcZuC6xMoGjNE83ZC7b3FeeasQl72kv6d5zzkR07O
ebS+owml0c5hmC/m+fhWnov4iN/biAe7rueAZgP8aEhZFCLNH6asBo35bBCq/VgXr4Por0NiuZWk
WnH4dn+qpETu07KWblG3CsabjRTZb4Cu+P4cC1rUJqvm2UrzowWgJJEwxGC7v+CQBED2gW/oTMRZ
ko1j7yQVC5KP4Fl/k0v6ZRUzYDgs++kL5g/t9EGB84khIPfNQpLB+vVsziIvmKhVqQmXAlz08xPE
0yqdAcVqa2vugiPfrdFvQrRESSyuZUw8cfFdE5K8velbW4FrjAYO5nAeBFqU8b7q9UgE2YDo+GNs
bYx0Zjx8COB3TW0f3fGLDGZ2HKzPhIJ8ViIzZFFSvlsGdBhbkDwB/HkVXHZJXWR2LGvtu6XRh/8T
1entKI3kJRtm+ZbFFmMrz0SZaXXSd6pp0VrjJgEcj4mWw85HhBY5yJPuh5Pii+k6PovvxLmFz5ng
DMM3jTxcWnnV6+/NdhsJZKsqFB0GYUwiPYDXv1yxlVXETrJ+IYZlWjcjl6w1dV9FUzUVz+A39qMD
hr6e1yo3mHuqbuAU8pE4HAAHopMJiygbgTvnN/0mY4dQPz0/Yi9ahI94Ukwsrx2C14vlyiNl2uWA
wiuW1vhWwPBY212fZeI/o904w1/mXEjN6YMLfIZNTpjNOqtdYU1VxhG8Et83rVm0E0E4pGwooucU
YhjyFlBeP9CFCLRSorboqgSGRZz99Mu8upF+4YhxKz1MhnO8BiRiPGQC3veHYZjEG3lWK/ceiek2
botvynAUJNiq6Se2sQhfC9Co/13VPETsamsWG6e36A3OBbhjAkfWzdXXQbiD6t+ptIN+B41K5LUx
fY1IevE4BXFe1mbN8HPGNm/LjEajKyJLW+QJayU934h66pAN8NrSREraIfSrQSw4Jnk89kvjLjsa
uwHqM1vr7MjiQ5gNC9owiONz8zn4HWkbwFskt4O3fAQ91s1AGKL9PlyFP6DuCfUQf4Y6HUAj73eD
hH+ffIFdokIsHkh1SkyhZPWoPRLVhaKydb7cEhNQnEnvH/e0zCtUHQY41EibK9Dx0GOd47vgehQH
mSWSEuZMU11bBtlIbMeT8Msj99JZitSnPxeK41SfR8+OZ9sDBSFLLAjD7QgWcV9Vy0hvwuRwLMu/
Z5oeZl077yRmFlSTqACfRw08IxT5GwaX7XT56Tg6cm9me7HnMmlwkb5DsCs73XCe6TMDjD6ihLxd
munhxp+SguBHNsQNa6L2QBiUsCGYtvD+YDSe+nK2BnCILAJlvJwrZaIcnSAuIqHxLtejWIdcG3h6
QA6IcVmPgDIBMlMRnzYkVTYWap3gFaB57CP7zPHzZE6PWqg1w9Znf4wiwhAkm7ImYPTcu4jdznqR
rrbAHtB6HF2kDAcNMfaqk0nHEpOnsDFA5hjmV1ukmNYiFMZ77CgrQ48v3MNsP/yrRuBt4OnMl+L9
+5sFw3GrTb1VwoksOVOCujOfv8w3pa6Vn3194oGGWGYzBBfF8EQG0yuXX7BUxjbqMTxt3kgHfeaX
jqh21kGl0QkWkWbif7T5qxgl34AFjXjjHDzyJzMV3I5ooEnZC4CfrUAx8tA0BjmqLFW6IYAs2CXT
E2Jt4TecppE20ucLa3/1uj3Tu6kRNtsEgu9A54oIEvGcMcI5kufCF75N0La6fssN/AGm+vu3hHlQ
wf9Qjw1qCmlUYoaMmywj0afC4bX3xnxntZGJHII9DBdsMeeB9PNp2pBfNeBYp4G0N9/MY85WUP02
OjXAabby2TCghddY4pSNQQejNtWa+wk0khdKLykBC/cG6d+3UZx6w4/SeBm1M74CfyyfvHZYVstn
L/eA7OCbXFscpodwYp3czP531EK87afRCbsZjQXzA80TjAATBNIjphGF75H+/wNQLzvNUciogxIY
VIPgFWbbspNeO2tGvM3a/zW0LREPNo9k7+Nu7sVrx91Itzolty9a5xTa2Rt5Ihf54eGExZXC5cVR
LMoj3veXoJF/usycrio41v4wWfov8KDny7opwo9rq8Ab90Cx3xYxy0d5rxBojBtf2YG32LxDMvse
ftK2NVOslbXIxcnU97NAPpwJNBoNCgZbVDrSBVhJn9E6d7qMg7HKCzLACEvuM/cN6y65f5vEhvdN
Sb5nRpQTtHzqxpP4N1LNFaKnopjVf8Iggzvgu5dDuauAHVvl/pJ0kuc07Q7xdgwKShQe6Ku5TNQy
q7JZT1f2Lhu08tpJ7lP/vdsV9yNNG/iHSKxTcFKg5DWvaEbup9izWoKp/kLNGkQoAkAnio/e+c6J
bTMzcUTeL6bs19v15V+LdWgvcczIEutPGf6dhRNS+q5WMBcvu0dvKtZQFcwgV4EeTlBPJdFjJO4L
+q503ypzsoRCe+UEfghWh4ZwdIlR6+izDOoin2pntCJ4mQSbpEg41nEqk2Qz6xkQsbuAY94oVZan
aNlUmkV+8gHpflmG15JCZba0ZWL6Nz3N0QYpWF2YrxW8B0/UvztfNmlNs90ApfSMD6Fc0aykndeb
/jbuR6MmIXWV02gM6GWp5OvyDzivGJQRssYJed7Bl2QKt1Fc4Uqix8UH5jF3lvY80aiXvTd8zBqW
v8UCLC7nF1Xo3QGCzeMudP+AAfCMokPBcGbmgPmDH+TMqVRx5oih6/dvOhZ80mE/fYzUF9ofZBGc
iJ9dE4c258U/XTio3lO4kqHYwibNDY3pPRL4n9IR7KcZDFURjj0TcCPAmU7EpjDhfgPvLnRFJ0H0
v/N/99gui7uxRutj1+Y1oJDolwfjqXtiLppTTAQFcOVfvCSNUArSfI4vlDsyBRpnQyvNRu/qdLM6
yHDjDmoPtHWE6anPHGcegGyzDaFEHHEWOylm0FI8GQBSVR5BfpxsYPx9NJybt6gDZ/pc7CMmgdfQ
+EObU/Wf/yBqy/eqJsXhjhlIBz26YhIVbJYahX6YJZLjqTIg0xe6pi4q3Zib3+NkY7Pes+PCTGl6
tiT1vSYs8mrHwzr/UkkQiH5up/r9SZOQyJ8l0qaiubLZCcv+v/bLQi48js7pQi74RlnmMJtcIrHT
quX7Ag04qpNVERq07H8dlwVpq4CloeCOB3Wb9vVegrU3SK7y735Z8tB3vwVhguCc3or2UDPa//UO
iTgRkBfHahbCc7IacpWSDUxChTzi+y+VajRM74gq+3rT9hqSyVtmCpsokdIw6y1YogcHEzExDI5N
Gn3KRMDm58nMUgQswUBReoykwZHwjzdELbRiwflvHVOWWP4LT2YhMSk1SX/CBF87l/quhl8c7UUj
6iTarpV8oS1agb+LBz4xxAfEIwnxR6y1ZeH7svsZd/sf/MzQSeXWAnm/AnRxzlFzhBHEPh6OX8IN
z5EajOLZlzURTOTipvEKccwgwVN4yusrsDmZALAOxlWXF3MM3l/MFk528h9AxRSoq9msUCQBDrq1
z3/G6BuFY4oF8SNAgGBnvRwMDRGTzU5R7IfI/c5BhUK23gFEzE/iZUJZ6/srt1IUTDfndLSl+Yoy
XrSA5+wkAx+32xGdrCr9x00ZWncN5YSDGxHNsRbum1st7RipGXA8ees7p7ghcg1cY4IOUnwT4MMt
k8DCESfIx/pGWbodMEMgVEwsWdkEnZFsjbxhGa+wivZDJIIHbdXwnwr5wYIKDTMUuTZt0KOuLzqt
TNibkEObtvLem0bL7Ns8AF8e6g31p5AAeTKcbVWvnvImCac5xYQOVBgvu4GU2g+B8xJdmSLxz8c3
HdupSGrCqHQlbOrUg9katVQVXAEzHzmhLCdVt5N6l7mqRyH4T8nL5uIAvPUrSq6PCOF5QJ51cEEE
4qISe8C/oC1/vzAiig+RoP+EEX076j2JHGBrqHkwi3Vau+h/fYeqAlCVXnbRchsSH6/G7Bndt+wA
rL/EJxLGUvzf5raK1aqfow4vdZ2Q4yuLCa8qgv331DSJS2lJl4bZqn+4zbt02YThE80dBbwYLPF/
rY4IOGnS4AzNB0/AChCHP9AGyXh1HR4JpVPfnRSnrM5DfNFefT+o0eGfMLUhbSp/QN7alDD4YxIC
/xlsffB3M3R9eCAf9kUpBXOU+9VzHHwcHSGWkC02iWzN2G7jCeG3N3nTza1tf3loPNBKVDZVqvUR
ywLDRgR2n7CEt8sjxG3XRwf6p/PU/1ToH0weLtjKqyEsMTedNr2sgnQ8ybjFFiHffS/LxvflcDxs
kMJCvDRxR6/IyDHZd0gYwz+VqNUPaCG+jFeena2uCetanH+dsGGdg41TxBDLIpsMTI5GT5I/ncso
4adEVwzA1ocwLbvJVYER4yuxXIqCBWLNhiJfTUQZOtl8u8fxBD/tD6mUAB0LrByXrH31z3+0HcXa
09fx2gppAueO6t+JSaVZMhK+6lC3yrVekbCOyMxgirH/i3gcIIEpBuGoy/y6DD4I2M0Yp3oLKUB/
6RNITqs8NTAjIXYE2fkbyiUDxzkHqN3NgjlAgXjRkYJkB42jEeuIOzu4ou9gUp9wMXHe8v62rBMZ
EAaFykbWnMn8KtZ023c8IiUxlGGIvVvP6x0PMhQ7CvioYvVwA3klXu92KO1BcpWtLEOAM2TbqCQx
suM7ZCaH5OtfLFZVKAm1iOvG5iHMoyyQP6Asi8YZvEyCqOlUwb0+JSTpYAZvYp8GNmt9EVuV3F6f
LTiKLlnqvFPDBYcgZJCvbfaQeAALwIom8+YcSqrHmaBVp51Fis9BqRcr2zsLhI27wXaC+eev9Uv3
sp5wn+VH+0kWci1A4X8znPsq0vYJ81frEYl26Tx58cR5zHr3pXo4Z06nVZUCPIQuFxatvX2UHT/C
PCcaFCizN6/uTVAK/H6CFOxQRhfHKq2l75RS7Ao3Ub6F3hAk1kpmiIcl70NucqpeqZhx4c3jVqW/
0Hht3iNZ07xJfwc27U2TnQBajl7NdgHlbbLEc2ApHFTBZZ3MZVtJyptX6BlMg4ixsy4HWL8P+TTB
ZIKVc3jtAGy8XXrWB8q1ExUqUdFn7MEdwb8Ui2Tc/OQVzJm0HBkzF7If79YJRQH+x1cYXpDBxT8u
xgPEXu3cQIvcW0SvYkvGFZPFq4IDtUkLqq94VCx1X43f/hNjLl0WOVaijQz2Of87K2qXT2kxi85o
WQovKR0OT65q38XRUzyBwNWSROAV1CF/kIMgByeVEXQAuUA4UfcPp4CU3ZHNJuFilCz7cDL0uCeW
iSzYLKQsq1/B6jAmUGf6c8lPlLjwzT6rTx0rF+kVrYdFyfQJYshE5IHUgcPoke9QiyztO6xkq+Pz
MtoILU+DX5+MVlubQwyhlxjpzZC7TR94D8xo6KjI4pguSaYnRRLhpb5Tbqf49oGWxqBZfZpH2DdI
v4OOX5X2STdX+/+ClNhdtzUHP6k/4FaqGp1/RqhCSeC42Sfp99waMwUt5mlCwwiGp76XY5ehM2P+
l/xf2XVJsP2CgBekB0B82YA+zJzAGG7zbXat0GmeaXFmHvks0+e7ytpJMP0eF8Zo33r0afG5UYCI
htpBkYSNW2lrzmOXR2rvLQ9+6vwHCRBgT9xTb0XC+zwuqWirEahKuxaDDjBWS8b0JEV4if3+Xk27
f5yd9kh+ZLIg+eep8xyvfVhtsoNaYhZs9vnIFRdeiF9f7PGvdT+q2IK23/iqhpBo2Ukcl7b/37Kz
Jw0PVsz0UA7xxdltM/2QJm4A8fFtxcxX3ruLQKcN8pC+BtE5YHMqnhqF+n/A+EnL9Fc5f/JpRB4P
vPbqp5PM/MkbW2NUJsBns14qQ8nt73qvTlPuQdqRj6V9eyqxgEIUjTkClpFTkrB4BOWNTINy8LTc
To3PQOYi5Fywcn1lO1LB0YgUfDgOppoFsLfo/5TFvDL/1EN0zVRIYgGHTfh7u6Qn9nCKHjK9zI4m
cMarq2fI2hHHDRfhTncsJ2ZEO1F+RDfZMoC0QOe4OY9KiHfkm/h8NyYNPXzjVrMrwSyTc90uY2H2
9DfWLJgVIFyJ5HKRbWv4YgeAOWJd5jfLVUPuJfYIvS09oYKBZmqzBAhcCnGqxf9JHIvBDsrrKEzQ
gqIzQwWGZ3JZPBmULBpfg1CnnKaE99EnCODG6syARJBkKIRGS5/93uKSC8GO9667Y+ZZOAHIXDtl
mAVvi4dGWRcpNbtLz7v6EDs8ONzjkNxO54Av7Kp+fHfw0RO5hSPf/k8B0X9nKCIK/vsv/YUsTU2z
ZJNm3nZh1LMavaCcJUpyFVAY18C6mT2vvTr63jxXfMgtb8PXdSAHkEN3estnGB9Wjg6oK8JvN42D
PGkuRLEFqpO8M588+rsNsjLO8n2aikEyj5xtCUz0N1mLVSRPyM4TJmb6BvUQDwN9sBi4KOo2oydE
L/e1LrqOcF6P7bFcymjPo7lmLZaoBWyMQRFHZrdbV+ugtaSdt4RphVDfYN2iCOlRMcgGlKRsW7mX
QngBXH7pbxn3xjjIZOe09HVawYsMnjJzkcU07OlVVD4zh+JKEU9j6zDbT/BCnrPQ/SYRdNKMJg1G
TB8QsM1THbNcD6XXPcp0Zgglyi6We2TsDgJlBDDRSXmgKybCHAB6hHmIx40cSRzbYtnwjuFQFWDq
Qan2O/ofW7WD7tvR0U/07po5LswzgsDM/J689JUK1nUk2P4vYRufY5KMmAYI6ezCKacdNqkN2OxF
ev9R610UJbZN/PeYuFbQ+gDTuvEpJJ1yLqKXpWD3RO7OLzsRG1qGHjt6PgSTHrLmveM9XWouSjKz
8LvfSskHu6rZlCdzoSeVr0QRZwGZh6YCnf3uTIm0N/h7q1m8fkVlPZAEeN7QiWu10jPr2AZg9pzk
OIMCW2LHBC6i/WuVsGXuAm5u4AS7IKKWriabadlnGE8TWshSu2K35xx1PHeTBb6wyzN51DQCzFPU
f8et6DrkhigfHBtm8nVn1bTEowS2GzMeJ5t6hnJJ/XJ6ZThHDd5Io8oC+oTMiL1zqYe3cuodAsHa
MXEz7JYnDeKHQVTYC98zETa1Pt7M6kaFd37h6EgLuyKLcrGad8qbtUO7dkBmfse2P4uTlQBMsATD
oE4Q8aPIRbObtAbqCdyWiDUGuhlzR17cyibhZaT7lpK8FgZP3PODcscdUOi70PlgeoXWcdAnN/hD
BsTgBG2UY1CkRdn4PrP2vO8MqeQfs248saLxQ7Wg99bWOZaCl/FPAYOdUI+782VTHjGFkTgKILTb
lcNvcqal2ioIig5k4Bh/dulp1mVHRcr7UE1SvoW4Gm2jjUXMOUkR1tun9/iR6+DgOXCs+sjXSuOA
HxyBhS4TwKmAfdPsc3DVSOkKK1IizvFEwPK1bjEURXAz/BEi2WiJqnvpwKAhpwmTlL0z7HRxJycM
D7/TWdXQ0jj6Xee7cgH67B3t4dGwVpFPdNvPBzKdAF03u+oV0k3dIaYvZSL1afy+Nzhdm/WMewHo
05M1IPmNRwmnXov6T0OVNN/0cBw45E6Un+ZDf0zER5KgGmvjeWSVzbTAluRXzbVw4TNMoBpPmMKS
pGpmOsmdXtmDcfPfwGefOldipaYXDTM6lyRiVRiOdNWrahGpiMXQ8r+0fKpnl4BJ3ci50+IloxtY
lavTEtuzqWthi+uGyc14l78tfCxHhC3/pIkX8RJreN1L9xynWM/Y0FQ5eXKTifGruXdTJNgIFnwy
STo18riMDg+G8DFErT55QwJIA/N1IoGgi0uDhVQovDtaLABeUbxY8+nB/QjzYecnxrdzwbHEeuua
OaKAm/W3TQkKtliT+CpNGb+TcKCR5fPykzPdmLJMF+5TTACrWsBV1FMWtKf0CIqEY2Au4rkpZrKL
lCgI/BgCtdEU0llPtxgPcj6aOAn/Q8Kz6w4SbENI/ym/pBUaywztSZr4VEJ2q1+aKlnklT6vNfBy
TbXQSINpp4Fkg24aYiWrx4fbzD3cYUA0HbjhRsVGkJf1ZJet1MC8qCVQrIjMsxGocolnzxlFlrPp
u8iPciuGvlTHBf3BPZqlt8myHapqVBO6boayCYXPeDkhIBfDoWyWDYffEKeluVB1bjRRmZVtvzdL
LjC+Yp9aQhuZJB0+0ZECYN0ihvuZeuJfFIC16hiqi+9cZh9yjcjgnnfCup3Zyrbtxa7remVPtL/g
+xBJU82+mZ7xtVj8muQEzjTjBzlXV4dsMpiY3GRBqYxjLmNlronbb779sBd1Wlm8Ud52wXqJCZSy
k9bzJEjt7fuNo7ofVelmpWIV+TJD5Zo1ftw4t+kbAb+xk2uIEKjotFGGG2LQZ2gqug4e4A4UoM2C
H2HdO2sTNfDDrHvrVYqAuvdhPX0RT9Ez880U8UTn21EWs2mT4EZpFMvpjGmNu6y91JBVSyl50iRC
woc/XT4G4PTkgB1czmtuAnGuUQmUdtOLX1TIrNlZXIsOoyQXVsjvs6bSQqI3mcAP4mceqIbyjfpB
LC3VZ/y9YIAxFk1KgAFiETUoF18ECrjgVtFHbSd4p8E15h+rbEUzzJOfcAT2DL7KlIZoLAnrGM9Q
xnLYHt752i82BOn9QBfPYRzgxYu/zF2xGjLAAAgsC70hlgjoiILa++C6MfOicIXYbu6GTq1BKZMx
nzxr1T6gX3+wxotCqW3c4W2zbWOSffgl61k8uag28Er8762w2WTTzrtc+T3rCAgNygxMl/YD0Kns
amc3xQ7PjL0NJq6unQ6Z5i6z7aEqW4Ltk+wWC41tO0Vk21M/5RwqeYgjH3yiieqxmDlA8jM3pjmy
75kdZZaYO/QPWCZXQmw4/EiRGp+o44H6sm+8G15vk9mZrjiOGdWpsGBHekggK0eL+5IEFEkv8jQF
RaHWE/BeenSC5MlKtUZ8kDNdvxxyUabnVIc3XE9WMgjN1FnEsVIahX41OwWWvP1lM62GKtEIClzN
LlUN4PbQoCCKVOD0wV9DDZYaEHD+uQUX//27Bt84FcpKEMLKJ0PkmwY3G+932vtkR+9GI/+nVOWX
cGkRDJTbWP+i6KreIou8B7DehLNda0JcBikjjZjDbVwdLVAu0h0wV6ei9FAxbnUIGuVEXbWWbgjQ
fdglUAYYglfBUC1NaBLsNJR1KhahEgjcdJlEX9lS3rpyNFX2oQhkhJfjI5uFD4DsFyPzbmwG35W5
0RN2V1lhPg/Np9xZRbWgZQTBIhrmGb0pGwH/qqk02K6gGwMPeFicpTchEEAtT7kWCZwrmZ9Y11Q4
KfnQyyHwrcfNbQEUDSTfc2JTrmSfKwrFPbzW1Y+3aLyBiajXCDz6cD5qabcKU4rjCJxffyMDIjXr
oKVYWl1N7mqGrCsffMqQyX5jyNOgcGkPgdWNPOksapnLbAynZLhwRPeicnd8RMgCxKh+XGRO8FHe
Zh6Mvbbf0/bX6Yh0ktvnrwu9qeG7B9C4oT0je1YypJZUo8o1g2eoyAuGLsjeiPN8NEFrJ1hOd9Fi
qR6wJRkDRj8rkB0c0wlqTdKaw0bP3Q1OhlK8i7w319p7aYQlIHIAneEhG8k7Zl1vWnRodcvh6ko5
tqqlvbMVE3Ac+MRA5pZw1p2P+Ned43cvdkh2TsvERt7YN457AiyyeN+aCw4FTS7EIZP5cENZY8i/
asTycPrV7t+OuOWXzQOWw8pvbwa5IK/NlSnydPraC9La7eK6NXtHMQfvzsLorxqPU0MSM82Moiim
ByEdwooPBbPPzg9WeJ7APQkMZWrQr8bGHp2DGzcQUgC8dlwD4SrCccOeHolMkFh/YXenLOOqUrBC
R//KTK1B9asE1p6bZ7Mb4OfHRvyefzqd95a+7nmcs8I1m2Hm5F2/nMHe5cvEbs5jFEMt+/tc468Y
wxypuIGGj01oEB1sxwvIonOu6XbrIX6JW6gB67R6CMXJb1pAb2vlv6xga3Unw2kWEi4DNCzFyBRq
Tx+vX0crDQvNUI8YqkzayOToFhq/VEc1mrB/rBnqeJl0hTwrJtAa2ZKZ1SwMrL51SQQAoYlhQWl1
anTS6/t88uaI3v4bwJ9Gt1mCB7m1O/4GWofvDkxEYfcIOkbwrXuU++AS0Te8wrshceJipGjjXbnW
WcLWrR4oqgCZuXvBd1bi0LoFaPxtvhi/pohW2UvIm/11rXhA6zODCvd7ry3AwL32Jclj7qHuphIF
zzU51p7syMb00zU/4zRF6rLmsbYt6JgSTEHeicSaW803NP30QfPolnS5kDIPyevnnJE6hHLbxnAi
WOtCOIGRoSF3H0J00xTy01Q8su/CFW4VE8uBDs54RNmv8upcT1rYELMr6D+0LWIjOwRTYI4XL0qL
aPTVzyOApVvHZfuowT36fabaP6CtTXK6ULFXgPkGRR8NWD62xAfoVL1Mkj1PqKh/sJNJxNY+WS6S
NTvPNfbLt9STPDI1duFL6OIQiOM+ee4hMHJRV638+T+Op1Zfl38lcmopgE9+VP0kPlRp3xIDyZ8a
4k1Pgfvxtt+2k5BF1hbD+Zz7vlKypHyYdH4uWt55jLU/sjbUmhqF/hDXFLLzVqf9JAYPUk3GIhV6
6M0IzyXbgGaFjY0+yuI0Gm2coDTWtXdMuByi4nNzB2dyixG4Id3F3TYN0qre6ybIcohRrinJbcWn
mzdQMhhMJEmZdnaH27AbYwJ4t1CWUGf3FI9AtDDsQT7O69QyAvHp/HSQo9PEjXXPUkclPrY3SZkO
pYiEetKzApD1cv1FzFVoNwEHZQqYlVJ0fuSOHS/Cgc8E+JbU6uWZSY+tIWMDVSJzgro84MK4cB/3
hwxbUpWnzcxNuHf76yNnuVh5opISthx4DRioIQWdsujDaABcRDZypHa1BiOI/TohnPKHhJgD7SlP
ivMkapjdmaNsPn0fd1O6Mmmo53CnO019W7JcSd0mv1w2O4NYKzfafOFhkdsYNWsEBmhwysXrTaNw
11WGpTrHDepnWOaCtaa74GIHWFJKghA095+HuNFTXzoDxGEy0N9SH1WQGSnszCnQDQtKQotJETRg
UyUh1VJUoBLUrgPCSFgAGGPwVfVUTdwYGy1+2Ct+x/vml534jZ6Ui+/HHVN36oeLz9KMVHCnyk8r
snHk9k8tY3Ui+tAedcl2LdfUREVzhunKIDFuusRLZ+kf7amzZxnhPrCL4DOqfzoyTjkLGu0oDqBk
rlLHStNXr1+OueQmSa2rWelxGAtmhMhqHMTDW1/8bpErZaqEoj2V8w8Kb6Y6aMS5P5k9oKwhFNeU
R/zv+nYmXHFQ1y4hzkPBcewbrRdB2ORXNv0axiMzjmvFYOvmBCCrz+T2rdIlb+aw+YOlPSG5DOT4
rgnj5228qaPnRKIs0LbjLj+KD4wqI0bKj5sgxtKSRWgyl5riMo7kaYE9nUm3/oeF3juHJ1M6VRlL
1nodmAIyCYNyHZOl/CSgtx5F8pm57UGvffRwbnql5jBei41077QBXM2YtDvp23gegrGRIinr+/YI
lunI++byMt+MV6R+AYkDduk/csyhX6z5AB6vxXkf0P3Q/53e0P7l8MKVp9J9EKne3w7mymJgNbN5
4mCVBICK/wwwy31FpDhmwsd4CTQ2aFkcoqKfHAvfvQRXQCm/9VQGAc67Yv1VjoW5KKUHPh7b57oz
o1CrJXo301xbAoibKfXJsgNDmDF0g27KzHP7nTT65VXMHfaZKpb4txTDf/kh3bPsC5prnVfZUtK2
YbvjTbHHwznLTfS3Wey0kgqW1/BBy5v5Qfwx1Dhc55G+uAFu7K336DSdqfbt6997w8M5LM8GMMBT
geO8bwTH61sC8ZRjufNw+VP7wyO9/LhqDRZ0yKMrqcE8gioOWGHJ1qRnZXa0Wp9rFqE3PDCaYhRy
PL0RmkiTkCa3VieHQhJjQIS8JnfpsGaehdn6QjFyiEEFJcsWy+dbElHn0rB+Q9sSKtiESdt8uVrk
13chhFkCfab+WpsJkuUF/dmJKmfgjSLurzfsK2P6iPmSSVnrfBZakLJ/MMvjA9Un9vc5LiRs4hJ1
LaeWL1u9+BV4S2kZlsXeDyjmilED6gP9PPN4ulAj7aqTfyISwa7k6pdZhrdWF8yGoZuoxll/82Mx
MpIrwyGL7Bat1r3i0E0CngtorOuX40y+4MRFXIrtWlvXMsuSRmlHHShy3hcycEFIh6QbEit4Z6kT
5pGByPuvF7eNh4IlT1aVc7I/hZ75LBgZM/kPZ3uz7C7gWDCIIghYy3pcL7+LwTGmpZ8yy+Io2NOZ
fD82x3Ko/iHHyoGQh55RVVEM9dCba6RJ/w1jPVhIONxlqbyl81wD5mS0aDgkWiQR+biZtAzVGoBI
SL9fsXv9vj9lj+Wi2AhqXcpmfb56f0wHCQJ0vYCDnphbqkXQ/zBmqG6M5NkvfUtHezIZE/ho9i1C
xUaoQLOct9IIarGyx/r6FOfm1zKTzScZbx5su5i6FBX2qelXTk0QUjJXME1ekd7kDy7R59uGHtD4
BQSYWzWJtGSU0I7VT+XqI5tmy4aaJlDhFp8niVuD1K6xTVKBKq1KKQ7n4+Fhwf8xC4xnYvoNePFR
rUICyxH08aTCoqnoSCPVCf5ID7UzDrzZqJhwVdkbxCBWSl/4W55/ghprb4xWG6crhul3Dp0yrs9E
yhKYOhbg+W13cTPsqyvaE7WljEMCcrILkY6Qi7zmEBga/wT6gsSnc7WYLyUc6aazlE4QRp7iI0Nr
LMF5j1r7YKwiqazgyFbhwBl3gRNFSRsFrssBsspzMQ0koRRACI67zub0QVXJ73y20BJYie9E8uxU
4tS2+O5FZLMzqFjEnzm+qb0G8WzE+Ge2+GSapJpmTlBFN3vSy0b/fc0eyQvQQBtBk4JL+Q5sScx6
F/yjg68pyNZDtHxkkiwQ6J5u+ynPt4ooIQh++t6Z/1JJ2D7zF61crVN5TEMnyK7iO8my4QMjm2al
vKcR1IYTqDM37HQec41NKgxa7t6pLFowNkN3LyiptyDobIn57b6fOhwkC8HVR94ZSaYx02WEBIFh
ZdXmZ4lh9wcc1x2zM477mRFlo6FHjLZ6Y/fRluIv7qMOoLAnwSE0Kz1mE86rTbqDV1JoGdA5X3Me
B/qk2S6c74ZdHejAV7ktraoy0CTUkZSmZLvJHjlQQZ8f+Lq2IzAV2HEZxSQ5qZCpcMwvUp2rdQC5
u1lNNqrE5kpfuvjcUIUnVn4Ae5ekHFqbNYzKY8po8ey1MkA/lhBZ4VH+S2x1M8V+2SfCo4tFOtx9
//kMettSGVgSmk+RlrSrQGwGNDIUEaTFEvZgLFEQHrBnQiNd0rhT3zoB9FjYyb3p3S7C/1l0uzSe
DRoZ2c7jb7oTlmOSS5KiTiD8fQCzV8hZXAwE9fq3thPzUJV7J9XBZ0S+OMOmzGkXAQRLP2A3QwkA
8QIR3h3/QGqpdKck5cTWmxebEiQQcotqSDHTzqBkP+BEpRA7+lgkt7Olr4PVPIj/TybEFk+ANuOD
mPX52lZZzei5wNayzfcz9PYgiMYk6YWHeUAFIE9bY1bHuL0M44ELrr++kOmC9JKBisd78nSpAzd/
844e/+/TDZ9DTaCM7MHSSNwhtYamdGyLhsQnsvFJdIyp1A2g7wmsYKGu42iCrICKl/z3nb51i/Pb
MEm7bJmn6AiOpSWDNIgumVf/0l5Gs+6JWJYCa4bZw10dM4HH4gAgO+JHt6OTz7kqqoC7IRXfguMZ
Iakb7vLj8XSwSQeXEVKYnb796MV2h7ujsNE2wZHXdlLR5x/FVKu9WwwSRfEBXI3+0fWhMD67AFsz
g4zu6yAipn5T9GjN1gC4heCHUlY3tJTzYfGS4F0R59zaD4yXFIsF9ewJwf0TodHs/NptSR4+RVH2
T5g14qmZTk3Jjdv9THldLtwY5etYMNvGtwkJv7YKZxc7/sf/ufINqO7o1zo6Gpjxdp/FtqCPcdZT
oZrpqT2ZLcnAz1VWTeEQt8jmXzahwWc6RDl44RapbT3JGsukx05Kr+y0ChJiyu4KPQGCn7eO1J0s
A0sUohlZk3wZ1PN9fqJL0FTjeejojRDrLyUAhoHswZ0hL2tQTe09KPxzPEpEIyALJn7WAlNyOlXX
sAXoOFQ1oD7kky3rJdJVVvnzceb/VIlx9VyGP925YHfag24qMPWXFtd+86yrUdT89EhT9sb/o4zS
WO9Jom+wSt23cuSVueAYvhkdMZWM/lXk1dl6bELuzliX+EccNtsApNxsIt2oTip2novTJxCQwP+T
Py7H/XB+4EoFIbFe0Jg5tRATizFPOo0Jfb3ea5QB1DHLja/6eNj1lw/Xkk77Jt9QpA/H3jKAa1Gy
09QrsWEfh0J8x21WEMraN040YpsU9lULrw5sJP4CouLaT2wGgJxNk4mzwy3Jclg0Ht5uPTd1EF/M
ZAZau13scSsliRBVonyvXgGylhCmeMSXfwqBVPJ8+l+Sgm6RLmzj8li5VhQOpIdgMYVBbSKVcbbC
Y0onJayk+nSbGb4VBTwydKo+2sR+WA9H+vE8Uea8f0hC+TWS443wBQL9zmtifGyuVapufeni9QG3
l5jWzr05pB9sn7n5x4EgT4qV2XzL5D9hzR6dd2LeXta6La7NF6u7Fzt8c0VBQC8TPEAa231jAl7F
98E2b4Cx4V09L8SQJ5uhvbj2uqpGBWCla8konMz1PN5hXt0KA+U9i9jSZNKoLz15jeoABn3eFglc
/w0fSCqN/NIBPI0OEnpYKHzHUneqWvEnGF7+/SUkhBL1fd8U7LvO4dr4VH3g+T6B+hTq04yDi6WA
RkvD7v5WxlfZ+wOPRm8yfWJkouP5ZjcbHdVpbpNhYkAp6w4JWBAGLZ8cXzlEdxUMNDuR8NDKOVij
dR3pt/CHtHdghBzk4Tb25xD7NhwB+DHQkeTSkYMRzL793hqbt+rl+zTRb00t5JJTS7q4+ySkHV+R
eLyZsbqOEF+TpT4ZzadTeJ2EKtBsnGj3zEqFgG+KQKm8ItummZCBDYnRIEcSQTWBLktgXLHo6EKk
oJn1qynV+qyDaVsQpfI+EfIlHU286AR0cUwDetaCsV4BEJVZbzlpFlDjFuNjjBrkOJtA8hTKoGBT
ka44tSJuryPUdbhswu4hYGatz2dcXiv7N6Pm+6apQkJso7xTJ6IMVF+owP1NH+uo/bQe4apyTQUE
wRaHQx+W0I16TA/314w+7RRTVxxv3cR3CSQVCJG9nECjzLpIhekmpSgJjSTZ/EyOA9uwte7zrt5e
tUFq0vCkuzCxfpWBah8qMbZZf2xGFgSxWpAbsmf+79WBjlCIxPRnpbcKeE7RiaLORcRHlViLQdKe
xpxTD0qvVsmy+5qsyZFcbRcyRg5OFiYS3RNqt09f+izzR8Iez7buZGfj7Oc28jeNXF7GYdjl32yw
zEYbUkHsCwteTHEREOWS3ly4gxBy7fEny5BZD3RVz6/iYgabaFsrh5ww0DmoiF6hvOIsVkXLjBZR
rNEg2Aw/DpC8380vuFA/OgG0QqDYRIU9ZL/icZppHH+xMbPpb767oiuDTMaENeoMBxxyhKkLFzJE
Q/pJc35cFPlp8ROq44xHsjSPU+Ku6V4PbS43bGg5NXJVtmp7+6l/HDGrCpciN5gvuKzdnmaROAcT
rc7nx3pxn59gSMj8jZLIpCnZtAvB5PawQ9kMFrcDiZ2UTkMcBeLW191WAvAq50WrCKu1SYU2bT+/
+rte5YvgCjdgCC5N4GbxNAtRPFJgXtF+1shVU2BfV/TQUyGOSF8ciKs30LqC+r2tFgc2zbKTizwn
zC+/W5w9cU9ntZyN2ksdHKBNo5Xfb/FDiBqlEQDa10W29siLrpXuZ4hiAtf45AryRv36YXq+RktO
gXxniEjQdZ0IWKlyROR+U5yQTHNDDMTsE/VLRb5qheNEndZ+knjK44L/jfQzs3Yay7kpzKZcj6Xv
3sWriPN8TC7XRfZd26H0S3c73MUDwLzBXhNVdX+CBX/QBS3IruL3ecbg3T78h9DCW+tK9i3UVDzx
mjc6nFyPKmYeJ540FrU6BAd1wwOmIGvhen04g1MKCpI0kmAaRj7d/0KaD4Jeva4yt0AglpopXyLT
A+Vogsx8yAYMbxu6R7jY+dadDYF89BdPsucEosfwO2ZI/jfbWhD9OFHeV/8e2m1kbtoCY7vWlJqM
ycQlah+hfgfO0Nakl+4+775JL/1GnlhxRl0DuPOE3qALHZ7X3jJxR/7ySf7QHqIuv8iyHycBakd3
UBKSofuB/yg8So5vBvUtXHtUmAZ+obu6yaMhR/VUQNVhBVK3asYB1qHBszZ+9cviPwp0DQujQhYG
yfEauL73+Wh6QE259pD+Xn5xym9OQbMIc2ikWPbsdgPE1b3JpHEzkXvXJiPxKYjBojHMjcn+MJ/w
zPRTnqDLhc8yn2fkEvsjo2ohcIcIMRWK20PBgd5qKPQ+P7xuGOUzhzlTkbwI3Y3l7N2ed4/vsLrm
I4pNZScJ8rB0Zs0TS5VZoPiPRQjrgl5/yk432donRs/7mbZR3xHTiZfPT85VyY3ljbX689KZBKPx
t/QGvRxeOJCkbCGKr5x0/chXPcaUNDOyJILr0bXvPQ9K0KNChOoHLIqG96yHcJkkY0U3JTYNfx3i
sEYpbj4iJ0kd7XZ69rKgCI1AnX8+evCS3fU4mspT9SBmX7hd4CXB/f/WDvnUdYAhBgqiKwICgVvS
t0gGqVC3y4S3fI8UDRhoyfIYZNLZrnzSzh+vOY7hBxh29fxLOT2kAVgJ1LBLco5wlfYl7PcFRTc0
U8jrrGof5jduHnqbyWFe/q9b6NbcLLQa6VFjVqUwQdgeGdUnCYmh7c2ItJxitwZ6LhAi6eUCMOXt
h4bOmmQ9owpOYGv/ZWOnojJLRWWMKcf3+zq6/bb15mJdNfrLmLtZmhDbBvDoacNdYShTTcgj66ls
7ySxWJYQOz2ZnETz1SjwG1bDNmNEz7sb0v5mqCCnuFWWex4w9Ki1XLwj1zLxvYdLYYjK2q5jnVAh
5aBoo/zbVC9cR0H+npAtgUhkJ044ALPCCg8gNoQvL+4eevHHNzOIMrZy6NlRAKmYJrn3/RYFp94b
+I2jVbXDdhh/aflxH5aTtpncrebL2UiDFXWmLDSr9CdbC8jiGv9gEAndyJkNX0CnluxyFzR4tayN
G5CtyL96JbJHgz8Q5h71xBKESsMEnE9nlp7p1yFrqUXoCu+fdhGMjlLm/Q4q/WXkVAjqO9+vSbVV
oLyxPXOxM0sqKVFKEbAc6+/05Q2hO0MwinVuAfp329bidJwo+rOvT/dr1xHOXYYHjDgN+2mr0VF3
OHw7mT9R+tztkcF+R/toFWaKuBIHLDc3x81PZAFs8QF6SV4TCaP1WXCQnkNoRS0uv9lqMUJUEG2l
kqo+CQj6/4MH2hiAAFT9A6DJegEbmzcgRPBznh3lVGzHOi2+djdlO1bGJLhKR0xMRw/ExcIfcLlj
qKzmRg8S3a6DJskHB6/FsEoMeFXkbd2H9YKPGW3c/yPSNtENSea9tZBGbsrbBNgshr9ucKl6WqpF
ynwzrtrUMk5uqT+rBnKeRfC18stLAQTcHnRTxnv88Zyq+gVIEw7Tu65IwVHK5ufO/Vp92sYXSu19
v9wNkASS+UQCLexIylucIFlktNoTrY4A1yWcpGNJmxbLPyJziNDzTCYKOyogO7MKCNN3+agJELOf
v7cRdobTpnekvaBxZZV7SbjEvRKt20rWyf0+ByjnykC/LIXwDjxG+0JVNIP3s2hPbTD7iu5ve4x/
UWIs7Kyg8JIUOFSbjaXGyUl8MNUmr+FGh/IDe/JMh9joDZj6j67idcBMiReSle3JhEzfGs1J0V1W
Smm9HmXJhEoYoe/oNKq6E2hA00Z5kCdk0YI6j4IWmRorSPpAOeoNhCbMNsZKT8FK/esixjB9ulih
Okyq3wwPlHxzRJg8Y8+J+uUujWoasXZnZzAYVyQdJqVm8VnP1GA6/aqadTmI67LH0Vq1W9uFjr7e
bgj8jm3hiufFaS08UP46KmuGh6ohKK56K71uhWXmeJvKoImwWXawZZceY59yeHPYpownNDuZf0Ip
S6XeTgBpHY6ZcoHR4LZr5nbPWCSf9J3+zSXDpSJVLzKdsLg0ITInngkbmJV0xGuBlB6+xIYRWAG1
d5E2ZPqoAx0EOxgvPDuSz9eshJPtzj5PNw/8ctXIFY6EjDFX5iYZGmmEn8InC6FhcGmEg5vNKWNJ
+9rD52FPvDcyQUQQVilQkpX3hK7FIzkjI3dSgjL+Ev8HelystEcEfzqM8mvG+ZTP2pund4Lt30Wi
1peUqHeg8g9c2lFrlUFndN8IS73gpagkf6lLBg82WOiqi6Hlza5vLrwDMW6IlLGAjQF//6klTvPg
LZ62gV2qFRNgZ5qFU8kCjtKLkR3tiu0rZ6Vb0HtrDrqZMrsB3THxoBktlF/QrYYnX/dYzwZLg39F
Qkr2+lOM90fIOxignhjDVEkTc+UfBY0KyUBPc7gMHNF7uBxSHMm4JJuBllOg68JGxxy493bkf/11
/m96Kf1gnebYkyV0z7b7Ecz1gEyPcPxuJOQhoOttRN5xLC3ex7MEPOL1RbtcWBaxYclWEzdqxpeY
qGiSuEkhuouc2/CfRjrLTIiDSyx0PK4IjjszEWM3iIxq0NTMmgXiKOFt8mCcTL7NAV37+h3zS1EE
LejkevUc3KL4MsXSBch0de6qveBXzKFh/86p/Xk4Q4YV7PibCqON166IKdGyhwvqfmwSoBgiAL1Q
yMgKuTmgZ7+KgKiXCjPHrGoA7iRnNuAT7dDyx5wBjLqSF08XrEOUysxVc/+ZqyonS0vv17gdMOYU
5BjNs/YHfb6BE0D417pRVTUvcd3/Vhz/xxl02h9qyuSrRBJdRBEFCBONJmxWjmm0nkr3C7DkKaVk
l527CfqHBgTdw3TGI82LuybShmBdjHPhp2n2cLM09jbqgX/kkant3CsTQ14qLB0k5FQGNdq0804c
ZPifunxkrUg+Wh/9NvKlhp2p05dE8kxilvf0CaF63KeVRl4PR/28JXkLsEi495RV6y6IOzFMPsoh
mci0kp5okg70YN1csH78IKAP02TtSuL+mtfo40HTJIouDzkK7bWu8EdPuEMJmLX+mhIkkbYoIfmY
o1Q7P1wT6RSohL7LRAbwKMYdc2j5tpr4CLOolO/ycBqcRSGPFOrPfmcN+yvuMCwWdEIc10EfLp50
oOgebvKT1R5gzfQFQWMhgN7DueyjCv2T2V7vWn0qVzurYob4+B4Q8STT/JJw6wZJIQei1uyfdbsG
ZnjQTekq8jn94g1DiLj4x3I/l/Hu6G7pzcqqPc0YDrch4N/CCk1byEk8Wyx+CPJti4POZAmOP9vT
vIxVxFOGzgdk6ekKwsOR6P8iW5dfkuc6Gj30Ur8nf8Bly/Gapv0WNTHSWVODiygjFXpTf5kBKsn0
MDuBgL/wSJg9N5SNI/rapEeejGyRK/b5DasTsCFl1PpjI07zwPTa54CCZYZC5/GvJZtdgE+ZILyV
mO+ynotDVVGBy0e+8PN/Kee0O9T0q+q3869ZUaqCmUokvBRGt6cSuMdJTzcAUCbQQyecVZ9qsye4
3Ustw44oStJSLl3qjgvS0Y2tCW16zC3YuqRDDlylhz06iPfLH5K9qu9tr9yWmYPdZxpEl+PRKewt
HcmIZIsbjhYc/W4vB82nc0uJdOCf9aOGH6QXBAVO5MbYcTb45m77IyY43Lxcu9bWFR7XMLiLxveJ
EhJIuGYZ+L2HsqaqLY02C8hypc9hhTk8Jy+0cjRvedN2pXkM/Od6y1MUf9U6JQw1gMCN1rJMLSLF
WMVVYLzvZtCFONL5THXdCJdMm45BlRqd0ISqt7IkWlt0L+moyAY/VX0if8D2VrDFZM7ZDiBZrHYB
s5MHcyKRJxAoqUyC5XZGqJzWJM8/ajr8Z4SfQGFYwfGk565rBVHrW+FdaQAA2XQHjs/mwDeZC+Dk
2ZrVebkcPVGcHbUyLdGdrqtcc6A1EmiU0hJGzRrIbX2TPzbAMvuVf05oQsFSXXeTUEvMS9kxXE/V
Q8S8FUBTLoFs93U4HHxRUwhC+Lo6I9OK3khEIy6BNuxHJ4xWDut3GjZPx1HPGWJdhpbqVM6sXiVQ
61ohHkrhkTW35JjpNlfhtPJ3M7k67fNfTv/E/+CzQSiNdWW2vqk1G76y1i/JCsGVla+h84UkN3iS
ZdQJlkrAnAK29JzmdTy2j9fkM5f16Me7W7zEKo9vJUCjvJDaTUyTvd00sKlXWMv8nlSrnbK6fshR
KQrE9Kr7zQXfvH7u3hgsILybEhTSTmo6AcSOS0GTQFCbqtBoDJby0vL72hhJSL/XUSxcEWTwIpru
NrdKWAJRbdi/Hcy168l4XQzCRWe21mrNhymQ4x0c7yPzbZ3EGG5ZFGUb8v+DSqDKH/1EPq/CzGh7
ns0O7jerUXEannvWDUB8Y8US80U/86HNhJmtNqSK8SnocdtmFJh4cBJxd7Rb83teEbZ9//vBrVDE
GUglZSTj7YnFf5xGwQdtRlmXZKCFkjSqk4Yieu/gJ9cprt7STxjc5gbppLMRrhsVK589C3ynLszH
LE7n844SOlSkaHZWy+nknDYmMb9IEOT8nH02w6A3JBaFo3zlAliCxfT6poO59/DmZrdjdvTrzFNe
Is6s4RvyyqMC744qdovAhKwxl/34it6JU47xB0kNQdzAiJ0sRpyHDxVOB/pPHS5DjpmnpyB75pEj
9RRwoNMZtmEfQGgThMGcrdJOij1Z9lO0Gs8br33Gzoqzito7vMopwXCoIww/SabXLrIEibQ/sCwF
1fWm8aslV9qKqyqKbBODiCXZfNty/KjS5g2h4ofMCQlzJzbmdt0pSLqdEZLPiynrN8/IklUzZzwC
JKxFD6mVVlVPIlXLPsua4CURB2T1mpZrOfbOTrf4yiRS7bYg2QMDbMyeJF1BI04NkTI85NUE60jd
V16D0x6E+crM086CThZNo75AA+y2Fq4Obk4hDIyAmhmK5Whr5VDv1rL4X06dS8XZNRyuR3RSpI7d
+nrXt1UCxLEYIspOpTvLeeeZ5SsXofHieqzA/VZ/QukAJQLQUL64MBLsyP29NJeWWe4zApYMUg1Y
oewcT+qwRLaTXA2YEsF06xxF4TTedUm4BR9MbIqhUt3nDw1O0ANV04vwGgGvtFvzCNQXhMpA0/ZL
Uz6r4PHBtKMAQC4XZjtMEC4v/gYrl2bYNDXzRjXiEHcRJ3EbqWGWas+C0kVNaq3tZMcDQT7RJGHH
XUFZFAWyP0lZa4m57T19zAeqQ3eD3ANHlUJA0G8dGtAAIh4KN2PEzqziAAiyLkC77o0c43WF6Xci
fqzTOtKu/Y/T59Z/8XKt7dhO43mz/BnczbRTObZnwkKPHUEB938cO1m+8UH7bBlbSe17SP9PWTEa
lkfCYTcoSR6FVMaT1IZ2LcdOUX7qtiuMNV2iF0xsngkQ31EY3pV+Zm5UcNgGBX5Bw7TiFYb1FneB
MXCOWObHQm4m71xOfB9KbehB+1NX7ArtY5w6J0MIBqVZGFej2CG+9B2fZGGnLRUcCYrEYaD/IOVQ
ht6GV58BaYfp0YG2FGtm4FgSlESH2+aq7dggv6z15lioUFjFDVU8MaTmPXIduI27CfhmicQrMlmA
CRgEZiJT6RAdTi+OK9URYbfKhzqEyRJHJxv4xMjiZKg0SXs6krLmNSHNWNzsc1be3RAA17FmiijI
dvOlipntIwrz3xDQSQ0bdC6gAz9qIAu9bNUgCP66r4DdOpEsm2xCQRR/EYYw59ZUie5WE2WzHtFO
D/DOqrScRabh6eMFeNfTnvBn0IjDOiUkO5v+/LAUzNmqM3cl937TWmO1WWNcNdgOPGjTbwjn448u
nFfd9B46cOvq+kKgptlkLCKbmACcsiqxFD/DflLwd4VrT3U3dcQwmAByxWp/RMGQoaWxbWy85mBx
/MB24SIAh41dbZKxkCcvitOZjcX6K1hqChzgNmEEwTPFoZ/SXvWk3Lh7HcxEYWfi6Ui0jBCk+l5A
AXuPikH7TSUnk2dbRSqvMaKoBz2uoRqor+MUkXP24tRWvWvgacoCHZIBexFhA0k1HCBtC6bUeWiN
1rE2eM5wL4Ss+s5t4Ts4w8DdexK62zI6juGYQ4z+0hXypNKx7y8UkEYE0PUkbJQzwdo0SM0ySe4O
wzSaifY9Nbf3+U0BLCm4zADfHPCDkIqGy0R4hU4fQV5XXiw+8Gp+vzhdB1bpmJL0KLO5IXwd+2SD
6QUKvKpY8KiIc5GpBaJlz0mYUt3O8xUI+VHlzFWjno02T4ryj3nzb7NRukrF7mEkM066ctS5LCUs
tiaxsU8fbniT++YTb1/zzzLyqE07aLvitZLa93wgArfFyMfrmvWejlYGmoFEBk0KPm0Nc3ifvThM
v7K6fJLx2r7JDs1oUhAWqI22E45uX7QegkLHCt28UqnW6iau8WdRauzVNuuIkhJybV8CmLZFqcSp
x6AP0Hw+ajGPn2/IqmmOiSp2ry/5BIh7DGQLluYfqmTdpTHFnqRevNZzTa+8+DczQOkpgGN6FEtM
eHMMRrwr52U+gjYZawKiwmKyyuf1s/y4FOEaPf8hlB6ze3kEA72ETk4et7rpvRp8zPa+Tv+aV17z
zmTAUad/0/m12tm0jFV+NnBbM3KblXBReMOzBOHA8+7ZO/bhirzuqWSLyMsryrbv3Ec555GqRAHn
cgfL9bOEyWPYhhqZpEzkB5oY3n63gDJ9f1eamHROkww6ChsZrLRsIY/I0vrkfEuRxR8uFM4JIUmw
mRRv9C8ZGtDfCYdDGbZ5/XYoHnucz8YPNAv9Tn2FHi3bLS/7etv7OvBqxMMP0FDfloaf5b1X9hrI
PObxlHmU/nn7/rlHMTMn23cv3yxGS7nUlp7Y1ymbodY9+Uiv8TWT2K50NgyXD4ik55Hs3ac1unzM
BkC73NG+6cdFrkRLF+t0MkAXBoD4G9lKSv0qs0jA4CCKShbdd6/yCEcA7Jb6dwVM17eCt2j2gn+u
4eInfSVrXxJwZ7mq1XtfvyFlkVh0VgXZ79YUHX9Ew1YM68ScUdYJvcCxMJCWPZ/o39oWL42fEXBp
W+Ulvh0yZ3ktvAypnAL/I6lEPUd4Q/fU0M5nf9bTN9WyhAOWizOo3TA3O0YOsIzf6OZJfNooD1PH
O2zL/frQapzeitvmD1C5nyTGNPjwVMU5+yW5tu9zdO2vum5UjtKzS+yVPZx2bdFydmV+kXCTgIC4
opbUpgVn2A/hld7nn0SyQ64dFWaJbEa4mKCVnKP1t1It2KF8naZ+HgTlJ1vJdMReoI+gyRJIzYwM
FqbnCrVm9m/yFNXTvblXOmhSDKC/ra6cuUFPAcRrcWPVhAFSOizFxO+unKalUWqu1RVjXazFXbw2
5iZpbpfX7qfRfFt5UsR7OxdZjkBfaWHVY0dAG+KsEl/SoriC1x+HpGxSxa2OGCDN1INdWojpInSk
RQETw2DRWH4ZAcVI42w/PQeWLaFG2s/B9Km0meCFEWlea83BlEvuolxeAZ2JcSRluWFdxQ2Gm4vQ
rvigzpt1hVV04/D+i5I4W86K3w9ryw0WhjO4CQpg1tknYHQXy25a4nofQLyIl1nCywQYm8dwLav+
2eGIO5C80DXNYHqlsDYHldwBeIGlXNJS+g+jOo4HjGqsk1CFRXN942eAEwbH2UD4HVAbDlU0qG+m
zh1dFokDei8PhV9y38LgFZWq+PaCWzJO5tarWSnlwOFxlH90VaXjqA2CTAdBo1PIR3MNs0ul8Bpp
TFzhFxKSqhfa2Q9aTi53VDvGxqQxUA3LkGrKO0w+K9uJFOhmbAP0zcsGvMQr9xtYFLYoZD2CJyHY
F+e65F2QtPkoAxKcAk9zVLCj9JzBtxPh5Pgnp8IDjsv+vPEd+T79ouTeryQ0dbMxBGtKwZ1blymL
Hud8bSRU/wmsvsHALqPOmcPiY8xEVQUBHxiC8ef/cUzS9aPQdJkVRqD1QW0VDtK5U38185leecB0
SnVr82MW1jUVIEh1MvS4vyZDyKDYjnB0IveVcvFEmiuMBxBbLjotLlrmge0lksgWejQdJERNXUw0
4QWraEg8NfY3501dt25GqBblKeNoq617cJLvyNikubKQax/LU/cMRqzXDJ//FrqHcnT0Fm1gfAI8
swjQL7kzm/HAhsBRNckaBcw+KMSXfFEMHhM0IHkoHRpDJ+5WfI2d+30svpry5EUkVqK31v4zBS+8
59rB78rpe88MR++E5twByBDm81HZ/qPVxDXcjKeXAZL1nLB4W6zICac/Vg9pC9qOLmol+Gn91JEs
nvpvnbw2KX8VGNw4YUiBbou24scfBYAp3fVsg/z29ui6RDUA7DM5doGpmIZbpnGwPcYr5zEC6iux
YTC7v0o2Zv8/VxGbw2HiDvk8vzhCK0Kok80ko6rqZUUvvo1GcWzkLxshwIMUDadiA3LTR9AvNfI9
wSdtiwcXFg25cbMFuy5DetQAE1rCIze58PkEFb4Lr2qdVYYA/FfObscxmDMfP3YkD8lb/BP6IviZ
al6PS75Qnz0S5uLs7FnU9dObOThalPxyLZ4STCUDSHY/LyqCzI1Z+88978AIRb9QoC9bxGU7ehX2
LPTDljTgtwawTE9UX2zDN3k42yKVB7CBkXEbMCCcah2qvrOZVKL43iyhfLHHoO+foxwYuD3pcWmG
XzIyKOhF92r4TF7ZbPhOr7RGndssuAQNiJ8gl21sm1IUu3fEhOz83YTXuKU9I8/vhE8pdTQb+Z8F
zWBx8xE+gfsPjIWl3252oHozrFMQNKN/+zd8rPIWiTDR2XcFWF5BmhcbFT9SLe6M7x9OLuot5xpr
1e41FugF0+rjmidMtNaF6GKWPqcnAs4AUsgI4k3a3c0ScmWLZGNULZaUvUt3Ud0JuEFWs4R6enpO
F/sc7s7OChbIf0K2OxEYLucRQfBtClA2KdlY0GK0yzrdc0P8s0el9nTPh5nIqeRohhN/LiobqFvj
d7HdOTWWvk/2iv3kOWkaX3BI8iyuzj6XtP5g4S2H8axzSFtqlPWEhMXDSyHsKxIqMHX9+3VPBJXL
5j8fK1t0KR3HOVeSOsFd92Anojv0Mq0XY+cfMbjsJXEk8RK3MLkYbpP9T1sztqanLlyAhUXmd3Fu
YhB4BCZRbC7lVj8AXHnrgdjy4LhPK/TSccLDIeDgULmOvKYXlskTaYebTPFDLC03ylLhABo/Bw4s
MXrsPc4mQuhJmXHctLaRBuZaTutLHdWvMr4SrXY6aH3BeK88zYRyjBolhhA+TCYS29KjD1LZYoQS
PdqLEz24dzhLty4Gyd8N8UyK4/2EIlmaD3jYokir/QAOObBtLln2Zk7vgb31M7Q7evYHva/QQO3N
ODfKZjMHOS/Qi1BkcOHSp9zbsbX+PQucZtT9HxC2/hlY6aBos9fp9qtX7bdSGKsvY3AxDqv2oWtl
S5yTH4GpxOx8qHmXUiwH6ngaAUhabbPM2VYkHW27pizv75tCnNeXThR8cR+9z9hU2+gIjM3JXK7x
x+dFviY2xtD/B8qNoH5lzMo78MkZFB4QVI09T1qlud8VunRQVbL0wBZcIw27aldSByL4BtXXctQp
lzvjCIMfd0xM/XvBnc1BM1XyU2icDG3NysANJFQGtefx3+gRUWT3FKIx4ndfgidSBNVD1yHQV1pI
ZDNKmkMR2rTiN8n2YxE8GYecb25f5a+AGHzUavCcrPCXYcSkySDK6aMr4l0rwlW4f6u/5Qe2y3JC
N5x9JwuvuAD26xKP7DUgC91rUzG7ZpWxegXJnx7GzfNZK1m8gE9awDlnh+kBzix9T/QttB4sexwm
XWgigYBcAaplQIbVA5crwJaO77wQmkv5mhSERSd0YOMAV5BRot5PVeoHjAGY6r/U9941xzpiRlsC
uJnoWA3KzXxzmXvnVB63KR5Qm4hy7l1Xv4GtYcdugSlrYRG3HkTT6Yg0WTlMDvUeB5g8alDK1Qk7
kNFSpGi1uWnMGdgRWIxNCaHKOdiMiXLpL1JmKTGA0bSkXchXihjKyRZmPCMjXAoVaMOwASiOBdi4
XHo31GNXpok7ouKd0CxStGRE5fgoQEwmx0r13Ib+ha7BKa4qsxEioGQ4Mxl3L7r09GH7a4w9H8do
5zd70gtneXpezS2CHSwK4GvsaRHEQ9sMSXh/DDWtyBg92FJ/wisk776D5gx41pVCy3qhyUTEk+wl
LxWnZPJn60yt3B/Q77I02T1PzSe0Sm90rZL1+y5SKfkGda6kLyd25X25HTVcrHR9nzZLMJWKV4t1
KNlgcYZ5mhTr/t8PUHf8fDF88wXQKcuQtCvlUisRr5mx/QYwjgdqZPFD5ABc/Xg4pHnZRdOzXAyb
pyGwtX+D/qTPWJgNObEuloaLKWiyprXYCOk3Guaaq8L7axi9w5eqBV03Ie925Tyh9tCJu1+vk/ci
q/y3fFUx0TKCHuO7DGRL+p6nLtMRMlmrsuLclnYTpprOe9UCMm80qxfFGL0LPFwB6Nm3UxHTNSeH
sEEFDa7vbU1/LATq07ddI3RhJfVcwmUdMlIeEn1YnoxqBj23/SXa2fzESMoM30o0EOzhzztrdsjC
zDIzlmQ6lO9QZr9IEvWW+wexqIvTd1/3zltP4anrAkoMLIfXnMFuylGhOeN7TOykbQXGbH1ddO79
aPGTSZAdT0Hcb+MYqaqMV6BkuAoF8QwJM5q4wi3Zw9ujbP7/F68ZGIwnAReTWIxb6b/aUBfoJaRh
Sb6nQAsQ6UybZmzFmdsOcdKV7Sd1H/xHI1bpxq3Bf4xRZ65VdxsS7vYvgTuSH9OGsVCi1NDmsGj+
/Ryy69kyLWvK3z0Kxt0z8jJVvgP1C+RkAmoLvMrhVbraaYcZpa5LOtfaiZWzp8ySO2D+d8JGbTZ8
QpeLGBZYJrxvsuw9KraJ53Pw106Fr/aCYZPlou8AolKBRGdJOHWWel59ODw3cBQ+woDzIKU6iVxx
KSNIhF6vJiN7tSlTeamvy79Phd8grNjlpsKv24BLSAMzn0p+O2Lori3BVft1Hz/F9V66J+GstMQB
9B/QTWFAOObPCPh1uKO/n1TWcjxZVoy92SiBbjuz7QK+nPQ5rrrw74bvQ7VflfxYzDJoKp4fimZk
Hsg0wRSWfcUwT6a3tU5qqo5/Gmti2dFVFAkCPLhphBHYJhCCbLobD7uFSOLHkRnSShN6AVbOGHUc
KTavE02XOdDr3nghHrDgdMmMVePs98pFLDpNPE6TBd40pFyhSNdVSrgfqJbZKQwPjtTqsQoRIzJi
pt9oRRaOPySCG6je0xdSg/mb78nGuLMbeqljLjocQK46fQ+6Mtc9yCm8SEq+AgCyimasYq732YIJ
+2y1K/SKip0XPHdfgtg9QBt4HFfpeyX+THyOBUmLarKPKaHEEurMYEa4HCnt5gcABYXhjZzFqth+
uoi+4RHIcHC7MaQ7k0u8Qm7jbt5Gx+JSc7OGr8nCfk7Py4VY1i4ZIr5hhMFCWwlXIwzqgmPT+9RR
18POl0gGj4ShWx+3rkZ4D/qJ7zwrsnCIZBaswR5knvF+Hq3EhkWnhjaKn4edRrgTPChYaBcQVEEQ
GRQKVdaYqOgnZsQUi7CxHWpFYG1Oh95ZLOI8G5e+fAJlzkwFwWzjZIfBDJ8eXG2j7eIGIOOtC41K
qaorRhbJm2W9dW82/SCCNmRStKMcPcRZVLvZp/WbJBlT65eZcjWBAu3gO3mqrE8DTBTWN60LTYD+
2Z4IYoDC0jSRITPuzi1h9pEp07H87pPN2VUCvByvjMDNlWvH69zLjqoKCmTzNuJXUHN8HBbUjlHT
Fsm/XMjXDrZJimhfksDfSRstjwDG4K0T2LKwzyodfHS1LwxELuVGsUFwU9K26iZWr40l/CqyX3xH
vwqgGsI7vVxJlZHI8E/PC7bhTSV7c3kjWjcfDjLRqfZ+BQ2giYr2Om0NMixeqs+S9E07pGEwgQkt
ff6NCYwUyxzSo3DHcUfYPRKSNcyLwfB3HfFhK4U/R86AUn5qa/U/hyswe5L/lb5Qlh+rO4ggssP/
rNRB7u4K0zpz7sT7pkLuqST3QnCeWowtcR2J0NJQLxMHzY3Kb2H3u7P5ZHNNx2jhdffOKDHnIAaS
8Kve9JMPo74FcnoggrdZNeVoaMsEPwRVbxbHw3Fg/XomyOcFPy/byMsSpBSdv61TPmsfEE/KC0uF
ijRHZZ8QJuXZ+F5oY5XaPLP3+jdpcxDE04DtdajLo0BKd4Ik9XaK2ePRw0sEqGlKyRRpf9gPF/Wd
/Qd7GrzyFtXG0eUDYd1EEOINxjznqnB3Uefjq4rosXVXGgPGMu9syE+MDH9GZIefsO1pJRmZzW/N
I1Z3kiF1Z6X39w0ujXAK3uAOzQgc5em+XO0iwRyXRvt0mtWiXHQ8mP+c2MpP+GJkKfJZdnP8tW7z
3WxAkKnEhJw85eMFx+moEiM9TQvT/wrJL8fJXj65QE0SLtQKnGJIObyrsriGN2jvDrykhMrAThs2
IlW9xRNkVTUdzABMVRBtaYgtFdIaouI7dncIugVG+4gZ3ZVenaar8qEUpz4RBNcCewulanCWs4Ca
teR5zzWlxh7wStFy4OmYvAJZ22gEIUgRwWlChOjUk+iscOWZ8bYMv1oWQUgjD0MddT18eIOvM8Zr
gx7OohyIPE6DbVFagoTuPM4/Ox4NrF8Qx/y9MEUm6yNdSdpco4ylRE8mPHNOE3YpWFNvd7fBlcyN
9OXGGLjimIfSJtV5Rc5qCoQ2qBHJv5/Zj4zF7Bfu7hqkhVVcHK6Lfw5bABW8U4NXfCj/WYpGxi6s
DlzD3MJhCUAa3ATrT0BD9KDmR+o3vMZPGV8aAdzrwBXTvUYuls5RXoSucVsRHgpoYDcNeQhA6Hlx
2Imm1qdw3oPsLRlMGDSbXfvkFPRvz6ctium6PvOimJ7RVYoDLfH+U3hzfhYXs5CNocFp9qa9yafg
xU2ECR35X6YLkN2WbQIkliu1iegrgkJ/65uSiVBFep5knGHcH5d2cpTlSJYHOzjQKhH+o74SCWfp
G0oG5IAIRGrFfaMBpLrFzH9woMP7lu3CjKhrj+TAMGmNXg/G/5mQ2O/MvRd1ThW3R34ZB637h82x
UWKTpLijYxrZQzySRx4oYasKMJwn0q3x3+TDrCqAq0UisW3TO8OKUaBQvqQmEnEiI1VGxRwU2blW
03Wis2hCL+X0OM+olPsUOKVc//A/T1Oym9COeyHcT3eFIWWv3u4DfLSKn6wH/TAK1QU70pKpa5sJ
Jwo3uckHIfCXsC68CZHTT9LIxqcTkDu5xOpPXjJHMRy1I1yAeNKkwTxGDu7Vt1AZlZK3lv9KPQvX
ZHrbtPMSnjdds2MAzK++3pnQ9rEzQFQh0PpicOoO80g6wEQFqGHp2Yz+WJmtIeLJXtrVoMTVw1Uk
5P1L0jpC8VCwwVYpx17XiV/V7HbTOBY37lkexXbExYFlo1mIWBfRZJnEdsQqcWWPV7B+enpp6euE
o0AyXI7ptz1mEHBWLcBGbpP6QjCxyF0PW2D+XwFVgtWs/PnqmIQmWmgpztLdSYHFvhkTTO/uRyZF
feAWE2SvkKMy5GSpRm4ETevep8HJRsBJnTmCyyJdHIUmuArsoT/GNzkH5apWEYyH77qA4UDFbAJn
ISTKbryydr4V/cb1dLPQqiBUB3WKNPzp3VaXTbnha0vCIQTnipXm73L35KOHNqXTdxGnXd/msJkt
JTzn+yfLaHCPr8quoTVjfgXQf3ASQdIBRT9FLwSB6+gKpPwBjiR6CBULzG/+kF+tmqC0yeqW3JXD
irarGXj0znjB/03tissgns6ToeCPHtCIC/qh84D4gQ3yi6137rFwFzsMOh4ZLtdOkdyYRx5WY+6H
DlPi7UvSLOyJOPozatwKFWpA3LWFkA7+DZn/5Dp0i7Y5Je+bqiKbElv6GCTjRjQVLmYg3OBeTSVM
zeqN7dHd/hlT46063GdDErBNf5Q4T2WW6ZdPT9BWYtV+Oh4Xaj8c3e6VSRhSg940Ua2xPIXOayMB
JHsOfVKxc+9y4h3nG513xYBxHCQrh4SvplGPjqJWOLbmbhQbPWauJmGjXL0qUyadZ00iu14+Iunk
BWrz4n9qijuQ0rBDb6f+cQ+z3FqwM/9TLW/L7SFyYiyTJRuU5kGH+C1LpHWQqiciAAJcQV6l6l6a
5D/BV4J2mxikRCU31al4WKMKu22Wp025FuJpJmRQLsRKn61OcHEEZDppA28TAUCzpL5eCl+NtfUG
VCevQpjKidXoGHPJZCgwZTcXyRgk3omWh9N4oXB5tBHEv2H2SBZwLgKKXwxyHsec6LZD+Hr2xC8Y
22OsMHvjKbYteiWb2cIQ2BXG2DumLmoQvm/odZNkAMPHgQu3HtPiog6LQSqBk/UiLpHEXHYIUnpx
BkAXyHMajXOkKOOC+PMfqExqLJQUCttUi42RYhN/duP0lhpKWUmxjqgDErmTnrM0j6Fj/3xRjAAL
KIC4kE2yGC6B3Wd6xjbSkPuopHOmlvaaBYKJGHNYVYiwF1qhgcUe3qgs3o+0nPQlYHOoYZ6PgX+h
jME7SsvhO7ly628BJ7C/0fP3pgt/OAseXVOrUWaqlzMhn5FyV47tBoZgdJQ+KwBs8Nrg8wcLbuu7
I8696wYsosbQuFikX9NnlZiyUZo7ApER2z4w38Spx3BRiCcVcYsI/Mf2O+bZckwCouJ2ODF2nm47
Y0Yfwpjpyf2M6JgDfURnEf1eU78Zhe8TlEtcPNcLIZeK09woCrUxthtwCioDAFa1aMe14ivkEd8K
r5BDAaw9SXKsNwQkdVUZqRblhdbT1dKuHvTdXLIVj+bf4VYvv+Jgw9HjtMoiHLjjQUe2nTEeOBio
q6WCER4wUXDydgrssBqyqcHYpgsiHV6KO6sG1ajRplYhI8EafwVg3P5cn9LFK/OFTGvUxTtpmkuj
+WHvuzHJYOO38pfSnb3Yk3TEFCPJdOZuqh1UvyQ2cyH0rqRBDqSjBIMBK3hZXdBpgRyYPT0lsx0L
gA0d2XXsRwgyGfiojUaN8twCYaKjApZ0lTU1ZhaABw1eE/3YNGGMvjzers0LHWbh3N50TqHM1iTo
63wNg1s19wUxiP46gXDHxCgqh9T5v9FkUvVOXr+cxAuxokXdrgAWFYN5+f/n82qunVUKb3OutmWM
lrCvDAos8C3FbTO4IHXdH5IcQcuyqstkSRzLHUl+AJYaoJfApJcEVauZDrW7evyWJFMjh0IgzBwT
PzLO/GM+LtzLZpRl2991f/GbxOp89k1kxtn+hzX+VV1iUIjuLajaTw+RkjBu/xAVTrWJVtteHhN9
97+HJwoUVF3y1fMXRCt6XAXPeu+lwKQX0T0SNLOydirx+uApvXEyySlE2f62awToSID+o0S+rkH5
7FJ5Qzhhf9G59R2vFaCeLR8wTMyaPvGFC5PSPaEfbcK7C8O/l/k5N46SEr6EsAtJeg4vW3JVHTjN
UOhY8oZiNewtwK7rkNF+14UO8fto33xJf5wHoLO4K3Hii7wfPV3KSRpDn97P0susk9lQdhNcIIAz
x+8CVZfujjFQkmLCW7CUbKlkRVIawK4nQpenbwdOGZN6yJAsjajNpkslHh0UdL0tY0TuRO9bjX8a
ePoD1DSs7Yjk2Dq8okQapZicSKKmHE5tHlvQx8y74OdGc8nbihmAdl13aH6LcccitkOWHtfnVDT5
eZBf5mL54qVD6ZEfXeI/BMwLkDFpmMvWFfhPl21S+V8YsrzrmP7vHsE8kS9RXM2KZPeFPzgG/AZ/
hD3Y7PoL4lbUTzEArTGBiRXJYiUYtWy9bhj4SWRe7mIzuiBlDvaPjHuWesdOg3DEEkDgDD/FFMV5
byQmqTvA6xqSxfQLiy53CTfejzNz32ZEiVmhkIM5LGagWQlzXmFuQ3HsnPdBLqUqxNo3eZNJ4bpQ
7BcRwAcq/3v2NS/KueOfOzxx9zgmCRGL5Af1FF+lE6xrGC7KWhCnw0nExUwCClJZD5R/MaEI7F1J
RJGjCR2d8gpAaPDr7j1al6Rmp5Z4QTY+9lWTnqt2osJ/56+MyuwzLXayTt5SVfrmNXqg7whFpRjp
kNPEcqUlLMaTgmLO7MfUXPPn6VI4vahKtfNi2F0XX9MwFdbfTkUtbDit9fwz6EbqTFaFl1Gie6Tl
qsO3d7xxKZ4ZGubiolWCovmX/cicWgEgUWxaQVpGTWk1JT4JmUeJi+sMIhg8mA3DP+s9L/xJOue7
/TfrPv0AJ2iSUdoy9r0GrGqxtkOxNskqc2Py0Cu/3gAWGnvpHVHkxqpkdoWi5QNTijQjF2cXbk4V
hSBzFH/ZEnKyTL3gKfiw/l3CcrpvD+/XOBquheM5w8OnM8+Idwxj2UK+mOKcS5FhcakjEUUE58ft
Pg6NLYJhbzhdwd/pmZlPrrZOHhmVLc5WUgnvlKHbD6EQZ+4QeXFG/W64HaQ1bf+xP3cMiOBed/jg
BiCErtHhNoFmPKrVUHO/2AjtDPcQtY9r8VPS/gc9leLKRJfVAc1MQD3+EoloQf++vqHzt900H5i0
iyMPNGIaS4KOYCZtXE4xjDNSHw45PxUYlyExyVtRUQ9njFd/az+gmnf0hULBbAuK8ZIJdoXLSMG+
WFWJbNA0OXwTL77e8CCNwLWqxHP7q2NAxXnpX4TrqVkqbd//nsS6ztA+4KenWEgnLHkYHSz/6YN1
oIOOlpkLESIOgzlDVE9ZC8gumR+qLQscDHzMsqjcQ0jvo2q/sspKEjeJrD0YNUiCW6KEI6YoY8ua
mlvODj8jpq+5xWPQkOw5NLGAiBFyFfoobaV/PVyKCM6afmcK9zhxPOpoiWiUzJ5HSlHNiE5AtcHN
aSYfpU0BrxsoUT6dnJPxop00qEwFtvOzXD6kuan89bNNSojO0b+vFrGl9g65eaQDCKCP4QpST56w
HFx9459nlq+OGhSJKa8jiYlg4ywGfu+mGYa5Bt2hgeVQrrErkAhMi3X311k8V8pAjwwW/fM4UAZS
mMKgPoGJtgVIKvp3PVlwrHQ0/EQwE/vawhMrtqmcQLnLEUtvIrNyk5gxUjA3Nj6IueuleA5jmUor
VayCd9gJo39vHgBGy2KuaVPpdZRIUe2AVynH+YDsqQPVU+Ma35q4meEQtaphTB+XACm3DLXHnuIo
YOTn2LdX3feG8gg3jelWYrIJHcJTdjxQl8FNNcMndmznzXVQ65/bQj07aiRFCSN1TqlDEq39CXPk
si8M6aTGiI78JP9Cg8Ked1KUnGN0xdU7N5ujcDfnc9ZgFvNhWfRfWaUPHyaXpL74we0cqkM7JoT0
AV7qEF6HNlTw5Qyqcp1Xv4/sNpJecflw4Vc1/9XvvPJMPjSrMl99urt1MJnNPAux1KgpE+tIeATh
DEmacWU1cW4j3o31RKMHDipJaEBCCsalKxJXwE+uJFbyxpf+cCvoIWVmybnJF2dP60lGHv0dJllE
TcgFhVUdHZywwiDpoFu8JgK4sGk/pRHc+BMDJlmI8dS5L0xo1IGd+C4sZCbXj/trmVnMAnTkBaor
f/DOMlpjIL2sCmXbBRL3K5a9lvF617uY7ApHgIOYxvujVmlev+0pkHPuL6ThCqKmmD5oFpBz/xk6
KxJHITVxNo0TNNeWiuVGQzJzqfxpkYeTSRTR22O2VW4WBaVdJ8GGnxBJCET6Cb5NeAkgRNpajxtA
KvDsV8OSzJjoealrUCC6+2i3iGtdflmUyqZwBfAOpKHL4QYQZBJhW9zfYp8555nqB9Joqt3zzJRM
JTksHxe2wqXxXbXPsYaORSAhM6A7XdT/bqKhfYTxmqrjLcRWskCbZA+v4nr0WRFqDptidgRl0NwH
g0K7zMBXSw4owjJv53P29ymAPQKGQodD8meMHJ0da4yEJwb4FG65vDoESm6i17k1JNDaU8GQeCZs
018KWviB3hOTEF50SVow5a4A0sTibHa1sXPtmU5b7ce/Wbsl+2ITOMDKafF1JVePHd6wepoL8so8
oyamcbZG+1M2ML02AILkshxJni76/Ik19NKz1RKqCW1oxKxmjM3Jl4loy/F2nPTtAJIlco76AjPc
In6P93PI1ochHRCOxRhO1F7rxy+prn5toYesUV8oM9wjcisSXK7bta0k5glkwaebdwIJPm1MEeeF
kjcNY2V91g8L65+kDyfOjBXiXa0Z0jmGxGg6EKna6BMbqCdbvELzcrc1wtJSy+JVnyUo0yZxPTIy
FNRdkjwz7HmcMYQdrEFv020BMsL7GNostNbeDYvcsJtlPD9/TiiWExa1fYf9zkqxcSN9z96iiBeE
vvKhxEuxVIKcjq9uAxfWMJeLGOALHSJH8HILPqKUFhTW9UoYifqogZ+BQV5VlWuDrLZTyAL8ALg5
zmrOkZzWaINfhw54klOHiwhKoJbe/KvG9+dl4i03ZXnEi8VbgxIIW08FG3Om5YXyD53dnUmx08oK
sSW5CbmfsGv6DHAOnezLvoGzKDBVNo+S/fwj44kN0Uey6+3DdP3Kmp+O8aRso6OjOQhmOljnuxJT
tl2Fhl3QwRSsxb6ZGvBytxbkzmh6WWUvnIkrFhf92jYm6AIDiJ1rBgSeewIUkK7Cz/qQ93klljBc
WxeYRddIC8Kj0KMCiG6zMQyDX+ZbJ706oIDks/7bX7THCXQVyWljWNe/F0EfcNrCZIAjoFMaQayJ
A0gDtRoQQv16T0LsMqCGKOtWQK7di9z2Xhzjf8ofCpRlF7wEP7vjn3VNm5jJFEWYx3oC6Pg61CGD
x3s5u/NZMFJP0n4k1lcmA0Rbc59prGOUxOfbeqFdm9GS2K9o11uV/nVBzPUI5pT6po3gUsEVFk6S
twMpr1wlkRw9pPjtHT664sQd24PZ0awPQ6z+dA4o4llA9wvPyk+TZxiVZq8WTflgoqz4aOlSJbGG
Xm+DIhHVfQuf5cLDQRKIsqEP7BnukjKFpzRQVF2O4n1DcLOCa4bO4S56DSAMoNXB+UkETem8qnzk
yHXR4yr2aLY8Zjxot38TOvd1jrfgRV5nqTfbJB6ddsTQe6nFMWBAusGnX5O9UT4spS0NUpDyPj+n
rM+HaNiOFGYLYURSX4QVb8p8o+izdL3CCt+IIlxVP8pjE1nCBSGey0yLGCmoG3zr3soQKAgwNjbW
Z4mlZji73ZSKJarEbLWLFI4uXawugNHom9t9y6qFL0Q1WBkSQTTRk/BnwSVuqA2S1YwUC4Ama3G+
PSDwjL0SK4aHbfo2hkgLC17OjAv1BafblG0P+CQroaD0xWOBF1EnYs2Cu4H1XkvRYNZrDgbjeFlw
7bBaEuIBKq4V3EVCVoOjaI7YfyqDnvx5dxD2u5MrpERx0sTyLKYfbFIctYonuBB8b4+JBdC0im4t
UoxIC+z8465YKjOi9uOSdBH5sTVprt2I2daU8s9Hy3bXMKiwz92Jh7gEbCVK5aZ5yNsnmMi/jfEx
9y/Y6WRDRIdo1cGKfcnZq3y3dqIgMN+z5n+ey3jG/ZTzxTB7FpkKAW0NwbWib2yOXyrmyBCCd8hP
I56aKqmONsCD79WxY9TFdZlyDe47eKNEpnc0HV1x74i/RRskugW1qbWsCYqBK5OS5gLRI9nnza5O
APQJeMoRDkK7+SqXz4kdjnv6jlbA+lVmDGOiLt3s0eQsb0JOzLN0FEtnPO5KQ5SM3KjGtQkdJiIA
rzheN9WqDkg04qgauUs8nkx1iIFM01UJgGnJOOM8xpO6woF/c+k8sP0nec7+QxN2RQQ3vvukxizr
QH5Li6vU2lO4AO8N28BIpl2Wyx2SYkt3sZmk+7prDAyaUG+KC0Rgeef9cYfVBdttpQDEPUSFHIVl
dKrbvSwFhShS3bdWImuuuLoqvtHoPPgLizLoLnpRn8g6cOVYyOwK9EcJzGsdRDGPF7cF3bk/DzAr
aSnOIkLo0aCPhau4Ba/yO71LEqRZsGB6CGCPgWL8fJqTiTrNT4Ipb2SgN1f/eMdNbZjAHdZwWMlN
GNK6FcjXKbxvteFE/CXg0oeuRqk3vM3yD/Casfkwo02Yknk/MFH5iAl2NG8kvPnQz1xYb2BhdApr
GBwEQ7rtNbfrOORgEWnwiplrR7iBwOFv4AZ+yWiuODPwuhQlxM6SQwyomxFIBYyeznsBli8EAHaU
zyAyP6OviGJvTOxScuCdnj17IpmZBkZtdBYxB6h+Wkbu0ogakAlbDgpopZjbls8VCMSchLZQTUdr
YSpX1rcAmKjTw1cndcM4kW7ffT9fpQc2OKvA0JPiqsiRAyOWeg/81lFG8ok/AukD8yAgMSC7h1Vo
JQJbqptW+5hYSyMJBIpShHikLgR7bTo3G6XsDPAf9y9qQtltd+B4Y7+36xE/yRXUN83AXnoYm0mD
fOvjRULAzSo1SBI2UEbG2/5EtVsNLd1FE27s6LenE4Q4xCMNAfGzs4nxTQHeOjrpFxwNTVDvEUu/
ISkfvDK9K2s8yJIKEqoOuui9Nuf8ZmGdg3i0hFU45y/dCfwYoKuBI+UClqMl8f6ZUGQYcJ55Fs3d
wbIjA+uFZka3NwqGSiy4864MNOtfRLM5EaOpe5UgNEOiRmk21NwEIb+58ALejfVCrSFSXYCLY4By
XYxL+0IT3br5Ex7BrBPDcGIjyJInlduH9VJi30Cx7xk7IA9aIeDIXZr9W96dQsCFJr5l5nhjDfm5
yVZmFX+i1duLJ29EoV/eUi0UaFdUVeA2fhvmg0apW+1nKW9ZQFDPB8Hf8TnHqMEY/QqCOr0AETMw
o7jkcTBUDYFF5DrlD5IFajr10vzRkvDt/FBOkkOZPa3LOqQNPlDU+/MsESQmvQ7jdqR+3GRTBIpn
pp8sa9bE9u7WNHflJNc31KdOoyTJIG557yrkxgroVKFrGv5Mx8sCR+xQMOnC3lkYwqLVAqlqj17B
nyIHKYEDVNumxCne2WyyoHOBWwvhYST2FykO5HNmKXZPBKv0/2usvB7jfZaWktO5dJ4yJsgmtnlR
gSqUtZisLNCVeFfUOGjf+C4P6glJk7CtHzp4FzySmM/Vf7ZcyPDvzO3ayDmSZyXwuVq/FeiBvO+q
HUItdzT0gG4z11pXPj75naOyHpiiV28ON30VXrZ8nLsTKGY99ilmxOg0Bwrxhh10xK555CJ7sjsu
HWQLF8pBQXrWOsSYO2GZiMkvewAneDeQz8cxmvHp9ww6kcekzmlQhXLGvumB3uPt6A4Sv9dQdwqw
gho0KX7zbMyZoiqruT4gcxmk8d4y603jUckAi65wAQtTql551iimlmRKkyC8Eu8Q3UzEZoncWNoE
tWe1j8QUqfGUONPuBLfTwJ77DLSr7F3lGqih2flwotQCkmzd2pux0PG3+8i4BKoI0A8Mg0RDX+4C
lmcLCVc21V/ymibyZVuMJQyjrYuy02/v2jJREF7LWRzEEXTLekPohq4tYgjiFI6wRvBlSnyZ9gI6
wHa6CbkxxuJwyZXQ1JbzLwUDI4ZtUA+3gWkyIhRthsD91Kj/iRaAqXF+YDaJDLkAoCrqeq0ASVZ2
OJVKDsJvKhBEjnfuvv0Xw2qs+AkXOuQ31jhzrNG1Hzt8XYlUlu4LfSPOwUM5kZaj4/fXBNcoFu0j
etgTliEGdu/QQ8lPNbhq25SCvjWglkSIrgK9Q2ORDUG5zkiqYN2FbGPbktXjaedZKcapqSTpy0EP
SfQV1gBPkBFtiZblx3Xt3aqpdxwl71AaAEvGXopbDY2JudjtSM5gllvI0kgxZkaWfp7Qds0c71SY
lME7xqCEQxcWggmyQkkWQvI9ZpIS+uGYMH3iiVvtDZ1v2k1s/LNqXnMaSbDM26QkTmJpRojs+pOm
5GNg0DLx+GkqNCVo6xlmelZVrZtC8ewgHKcAEXeTZDdzUnpmkQb4IXKYPBERnZ/7aE/yQsX+6MYw
WiedwwOLOqYpWVelAgXz3s/oSOXtalCETYDOxeNKGN85dZlNa/5Cpyyr2EOxutzOrQ0Ummgwcsv9
UzwhDdqu0xSBkjRdenP4VPkVQLNjhZLmufp7y7zOUigeHQ+2k7ynItilMeyeHDPk6og1UGpdfLPI
ehXX3XWyIJTWc8LyuUJXC2gAuwi5yoRkgjyZ1gjSGIDgrVVNPWN2iIvcGfG3e/M5Acq+KBw0kGMa
uoe2P1uASD/iE+aEKxGvzPVq7dvMFCcSlWcnU22gUdSMDWI/i004lTyyDE+oUUE+EUUG1C4Ty29C
x9zST5IJu05xNDIFV29qexSYVIODmVcg9823XuvsJdMZWTuFGBn0QvF/7zJGYScBnAi8+3HxuxeN
wQTKyObxML/d5QpHInpKsHHAgZ7kZcEw90R6c+zlMqwSfhrVSqXzky82x7N2t7ggFh8JtGJUl68M
7G5csYDilr1TZdZJaajR0f3WrsdNyES12WQLQUWBZX2ZyGhvKqTDAuzAEGKZSXPwcokPQKtmNRrQ
3gsaR3vPG9jLm78mJdlduFf88CTcqaTOiCI6gK4sFNESYEFdCaubG8htmaJc44pUf0YHqjrvBf/i
iS1yVg9WcA0zHQLLBMg0oXrN4nuDc/yz71I9J2uY3AAalRzidVkPBk4zHncNNIlwLj9QMhw9sQjV
4/y8h1yNSB5mQEVtpKBNjah6UAsRzVe2uyE/H8vgnsf1GUHJ1fPH9exbn71SuNTzHqPOzpW4INRg
tWt/QLVcj77tVe0zxWbB1A/xK/1Y0Y2n+w9yGquhc5ZM0u5srs+NOoulGdewLtr+AgN1RQPljZfc
9zGpKq55IE5iqB2jmjIiCxaa+prroEI8HVhsRj9lGmySJnDJ+JguuyfT+mmSyxQGnXmRwfA8oCzA
DzaSDtRM9eaVCpvlustuT6CnP1i6v5x6XsfSTm/vtAlpI3LL21/ik1ufiTC8xgjVkp66b/HQAt5S
BJCzraITlNGBg6/e41nhd1uoc9xV5oQ6/b8HcV7ctCVLq5IRiftcuHDzIHPe4nUeNjTC5aDJ825h
EggLh+6aGbEghfe8iCrPb+HjLJh2/NXcqV+iURXyFGPvjLPYF3FAhSywd2u5Cuy+ooirhSkKVdQX
mU48tEKX0qNlNs4CSb7XThXeAAcxRX6bQ68l5w2S8WfwNdtYIaClCTjPgiUIvcrTrPwXwGlU3Pn5
UIOgPy6IK0/01/5wn0yKiOpxnSh4zyRYvn4iWBX+NjUMd8PJ9P3p4IhdrsjtwNPgpPQ7Ad8McyJj
rWgNjK+w2NpFhmxx+dOTIdgMgs7y0kMZZbNNIIHQZzn45Odbq139mbYOozpF8cdiY05D5kEpEHqS
sykeZQbrJEmiBJjlI8tVA5ij18Rk2+KquVe+KpJRZjYB2Zd0qbyI/fUFCR21vBknwP7dR/LpMj8r
L+cjvoB0l6qxY1FfwcFaEkQi5cMotBS6Xo0ncD4GABv7txeCDekgzcPX7dquDMrm52uUbMbJvAcI
sFzJ4ekENcevwpkwK6wWwOWkLg7ZD7tZTf36JXQ45ynX3UxcFCtE3bYs2tEL7EVgSfsjmRCpyRbS
DAjvOsBYvw4jf0fm2aQG0pSB3O61Xxwv1oBgV3Jxh4JUlWorwH65QVdEmvQ9oT9BVNh+UBnT1YS6
EHoOo+lRoiYMWuhSfSJxDAkx62mY4O5S1mOl/BIVydKdgp6YZwwQnVaC/oaCTC6C4US9CZPmRz+j
mxV32XGQPzo2z8DlH+ej0m4QjnQymi6SDg+R/2Gj86XfEF70lhJRTQX1Z5Y/RgCc73rL9nmKh45T
1N+WZb6mZkBzJshSpPvwpRYh5yc1gxrg8MSwEkZQ4YdiM865GvsVzrtakD/c5E4dB8K/a6uYDIFv
WkEQzTUj0tnV0nKgAV8eaSpJRQGzDpdFwX5geS0dSZMjsCQ49aMdloCgxG1gYcdrfXEcJhLTRrm3
Wf+SNhklVSn3w0+ojOB4q21eKTE2hVToO2GxRkCc6gxi2uy2JsQGaevnfn8NdKqpz7AYcz09gz43
eOU3W6K/zPlePAwprRy43uFPZA3IsHuGeAnjyMaJ4FfCbMHhpBGlARrlW+LeuK9p9+4WNohq52lK
f7PqzMBdHeFtuApQc5xUkOevat2uJtjsCYY24agbcqS4sADsSktAp89IJ4arCrd8wz6UeU1sadXS
QfzKUiAX7vo23ghXkYTNdoSzfUBJMpl85++m02/HCQKZiwhiJMg6+eSWcx74LlqPlwnzHEFef1FK
OCY6uaJaSUSNXZiP84CZAbfIxOXMtyRxKDHstCLRjm3D3r4Uh7tI5gwBSZ5ZSODX9eG0XrE54TfX
4qBU+Jrq3SEb1vFbykDanZ9GzYh8MyNZ354IrvzpKaSvZHqktOuM5o31VylH/mVCqfucwuaNeeNE
69kMrn8nmSQImgonRozUprqAIgVIEoPllvwNiMqj2VGzBHyvWim3iGYNRM2dGLH8HMvZzqOp/SkB
guObo5IhXC3aYmgFMMUYF43APyD/fC/sCoVvhz3lOa69lwacwsDYUMA9bcpZYlu7IGgztuJFNSOS
PFv9iU168UMYlqShFdxobCDrr8j9F4T7Br9wLOXMG1Rfdv7yLijrZyn+M2nUYLuRJxRAysAd5hvJ
kAlStTXykPgyfMq6bIMdBK2FGCzzgg8/9LyRzzQcwtcAAOmImQDQzBw//CYDO6/wkQYbUvxkef15
tbWlPKth1ZN+DZ0mCYH7bXtSg1Cdq4ihPzY9lmMpa3LT31iMQU/Ncm+7gGw/7xraVdIyAeVBqzIb
mjIf0vx9aLT5QDGH7+e4AKYb9WSUSMo7I5a/Z2TKUs9sH6kIQHYCLCR5RPF2NelzzH/3pP9FIbjD
IqWZJl6K5TBefCW4czCxMCKOqqLozPRcs732A/nUhENCLJfPCeIIBAFtv6kj9ks1ika0AbD2evrg
qNA9df8jBWKu8yndITz1UKLV6Nk17wsrgfRyhzw0VGARQHXJdIv164l/DGBe7OMfdaGizst59kBa
TICdC23LyXw+07CJdn/gYVT81IjyLzpcK8TVZHk3TWMIc3efurbECLd3z4L+Yaxtq8X1Ewu9D65X
zE3Ik6REnmdTr6CpUvfTWOJnQsytM0e2uyWKGiPDdEwXlQwRTqQxP7q8PS25cQOOYCCoBSdYBTvL
fUQKufvnX0BU37S4Z9Wyyuj0c0MRaOmasuWlI6AznsN9ZE8//Wyp3TD0Mqmy9OsKS/y0xmFg/M4W
VZbPXLJNC1pg3afT4goTTB425zqw8EHb/g/tRWH9lgQEz2389OIrDlzdV9cdx1g2f0JpuU0jQVmD
szfn3X2q35YLo7IqCX+aG9SoLI9syaXoi1I7WSq7oSFfJxKGbAbDu3dqXyeQPjSsrZ4GXZYn97VZ
2wdak8mHUmDzn2C73ZJuQO+xxESSVnAEZ8A6aIK2WCbcunGjvwCYwVdMmAZ6YIbLjvAmrrzFtaxC
MI6e4rP1a2f4MQf+PhD06fhDShmp+8EjrpD6fWIApcIY2T0Dng/vpyXLJeN92x3mQAbpRsjT3Ttx
ox8ydIh9By/ggvszuloXGncin6bA4Ujg8mYlAgJunfAY8iVEVw5J9RbUWL/suqdR7a7eQbLJci+E
iRPxkQk/xCJFnvcKXhv9zLVwCIrxX5cg5joym/F2+gGH1zpyf2ZbIHNk7iv+WhnGC5cWEiTQNcy7
wUv+E5oGjnGaLscxrAAesH5bavoHrBK5DDEADaK1AWK92pueom7WSpPHQLP0l0YjM0VJF7vouJ3A
U9H1OWiK2gChr7vdff9f0akUeBCuqEe6Jh6UbS0apUDIaqAUR358cKU22ngwsbYr+6P2IVWFlJ1J
oFEOGGUUjo5/WWC7Itr8vnZAPai/0unCmSTr9cT/sa3QCRy33qhjtPb8BUJysK+k1Mr3d/A5Vpxs
f9NHnAPaAqjNTKIKlhMlz6K7/9IITk48WZBKzB13ZkPAuMVs3Wt7mH4xsKgluUghTNrXt8JrLT5m
+3dmdskUCv0pkDtB45uUviv98c7aUZG6SkZDfih10yjMc5o2oVJKW9qcI/Tsacd6nfSjfCwDE8ke
TTQpVLcMC1V5U53DpRLh06zAD1WqrinCLUxpTiL0+iVUrRpxKu6cxoZNhF3SFgcbucKzkHKMlp73
ppj1rCvQt1STa7lIfQ48RsSTYAv2i2pvNeWl5FcwcxCufxid/pY4d8E4ZRvLKHgkS2asDIE+RWgw
CkGvFvRkO8O3wlPqysVVZWk0anSMRUphvzPYAyd5luq2IE72G1KXcMs7dt9XFLeIpatvcp26PzeW
lZEiB9zwYW+FCZvFQ79D62p7vmaCacH6H0WtVihQt748eP9UbUc2hSv5i5RmAcOVyfTSkv2oZYbV
8QsGrRVN3oxeH8ORtBKVZwIULY6CPQUrVZFs4u2l1zEWBrx/yg2ZCV68uev3tofU2QsQpdC7OOeA
eyUDb+Dljyht5Klru7M17w5w82MEk4aft8I2TEsKIjyTT/wpioMOHM+LKRFxVIpMucpY9ElwV1Oq
umb/5uZdyYwuRQRDD02+kW1upKmAf5XeZyXsgaDcp4IHEb3ntNDjs0avnB27uSlOIGdpwIon7tTk
GeDTyhX/OUsQTBDrN4ogqykvy9fhF6K6DUlD2r0uLm+uKLWPjh4zEgWlgTR9Sv+inCEUw7ewxe6b
Hngy/itIItqIpX8HUYmgiROXhTJpuvkj8/V6AZJWErq2wypibzBUX6xF4cEpcPXnoFu/oSH19S0R
A9PuBiPCcqTVtCOa28Ej6Ye40YOwcb7aYUFVDqBJNkd6e9SNqgxsDwqcz6uw/QbG5akhQGJpgO2N
4PPprwq4NcgNSIXxeV9C217CF+6mHctNv54iUQwDFhrMyp0VRf/X/FeTL9/Tf7J057y10omu/4le
GkmUIa/vRPw6iVP4hELlyVzu6VocWTk9x0oQOcIjTMy016PoG9Z6WdWRCwDoTp8jiAlfzBdS/+fa
kx4KHOgMxryYjB3b8W1iMENxJ7Tpve8Mgs3K+F8KhRtuHrOK8m3Z1Z8HFNOGIFYNp9c2tcCOzUX3
3iYGIKkbBY33jb1GgECogU7NPCCjyg0LA3B+UgRn3WJyAQ46ZzmUC69ludQK90aoJhw4ajzRTJF/
hnpwmUC7kAhYtXUtby71BA8aXSGpLG8nMsvo1tKyJzCYJXngWKGRAC8vll+hlK3qA4i9RViqc2zR
LcEgkbDSBlMm6kTx2MzO4/ZJ6+EYLV+u+ZJB6tzcw3+cB0faYPRogZePFfNV+UxlebEA0YxLHH/P
5CDoq+tP9flU9d+JuyJQPY92rrU8Q7KSOzw2sqQt0d3mDA3wbRalyRI54wVk6b5g37mm7iD8Raud
HIm0i7PD/oeX217PzdWoiI7kiB1seJINorIx+ZkcBHyCrpLRr7V0B/TiuRGUAlVMezRelEjpHCqE
msA/HXhg2HYC+6tdpuc+4xYg8k3+VzDeRiCK/dW+uB8SC1Gwy+28bQ1oyoOvopVRc/wX/+/lhGhM
2R74QQ/YtYgB/XjgoC1/9i0UNFz8+gX4zRaZmMMqpAqkthOav95kDECDf49yNlhIz6HuI5y1mJzr
3uamV9O1Snokt/yPhQc35xUHVH1tpO5qZkOBts1pRNR6DGRv5LNraExXf+48Rqk4S2ckYBl7nI35
ebSKz6hk2suVQsy1Kw9zVvTPEDW+niBCvrrlJV+bSNeVk0VaQCqTQKrRjFDzrLiJeHJWRLsdNq23
EqZq0SUy++oJ7GRezsyz8NoZ7DFhOSSn4kvs6F7wc/OXwDue11oDPB2OnniOZppzJa1Rqa1vghix
1CYDwM1ShniSTH4JdkkueAZ7PN6BMYyR4TCZKZb2iewDfsb+DwQbKHIZaRrOKs7gBCdyL0Ms/zr/
uoMBb4WrMqGxOtVuKUjDdp/ujgZ76/qK5Li52s0V4+zkZhLiWu/TgIBZZ8yHv6f6xPwlqk60NFDk
esDsoqh6wzIPtbSXCgT9LcBwi6cHAub8Eo6sMxvjMcf+TIdRNROq6kaloRU6igb25wJOJGwg82i2
DDei4X6cCCB9scn1oxPJRESx1o00HWpz08Zn15CRwd3G33r9SdTlqFfnayexTW5lcDTfbhyrqZot
kJ+hI71U6JqJFY3jfW3TaYvqjh6tiEGT4Se/E4sA7LdaWNGSDtzXjQtLGwSN76FdFGkkvcG2ioUe
ZUCC31AERQ3PxDsHkHzBRl27hwik0JAlSETxLG2GIlsHJ+Xc4jdSD0k5CczBaPF/8FkbFYQttHjA
W1DNeGbQKYVWpI39zvFvbB1or8nC4sYvGPdPy62nhO8cDrb9LEUIbVS5QbRCngVpz1FEy6MQoV/z
co3H2f0O/rmVP0R3QWr3XaRAYnBjDr/1Z81w3eoggZwRNJvke3rgcmxdbgkSEZC3D4zsWKwx41+T
6hYyIIMoRVKGiVvBcEYviW9wtQ2FlAz55GdiNgF0XF/FUy65GMLhfjbH9b5gzwgkkNA+Ty5qc9Gr
8c5cP+Q+4eXhDnKf8tET4j+iAJJ91WruTchhj/eX52+zcetP69a0D0ag+e7NrTUyQRtaTxJzOOe2
h1lETuTa8amDEOCr23eBEb7XAYve0L0T8WD8sbURhHfZ7cPLd8VNOFEVT28j0U6ZXhbOG2g4UkJm
mivoHVpnd2CwJLnwThzJ64krn47NQ4hfCTDLIohOYOsej91wSZDwbRZ6zGqckyedWR+6tZzhYsnG
Z68v3MK7Q4U+TzFi5+wYMVlA3mSzu/UP3zWtIOkOS3fAef3RFI02RAskhCl4VCWRutV4id/0cK/c
YKYciRMY403TQDi5Su/Rvo7s1dVrS1vmxswQxA4OnMzr0QEd9pn+W21+5VoMWI6YvK1RY3MRNhwS
SGXvAZ/ilTwve7whMM3+zfnPkry50QUCJrFJ9VdLmCcY+JH+zq4kMY5q+nIIu0uUUprh+czdqHrb
emQMOTeZRqN2OA4KzhSP0/dUZBwhEdxeZGIMQnpQxI4mO/E3trgim6ErPg9H916UlEMaAJhes1kk
/ADNum+9hCTSq1tCF+1OvkplZ6Jx/5Sz29CsFp8eONBg3maqlQ5YaMFmWDzmGQljLW0TgNc4e3Md
79Nce8b8SNNzAoDqb+fvHktzburQHNz78QOc8GGF95Bz+HGhhMReXwAyY+W9MOL6Qn54ljvxWzhJ
+dyMMVC94FmBShaiecJW/mw4BzRyIEK06B95lxdwPVgOGQWYdG9VN+CmCPS0GaL+lO8eSpi7jYT3
R5L1NS6VCQiINqlYTIG5aBFqvICQGh6nP45H4+Ww7phhShzMJmIuSt8kzRbvz+l+1J9JbXTTugz7
FzWD+eXJvgpO0ZrH1YTi7f3YPr76TDvulDncG4tB1FKKbslUomaEhNYfJ6lXY1WqFtxcVxaPTJ/q
GLSVfCVDITOTOZX3z4pCW7QAd+f2KTwBV4DDzvzvlxyZskMSyAIA3Y+doLQKxdwWe1v3R21mI83i
pXkbfDKbe2NnNXVR6dxXdZ7xXZ8JTbme5ICdbu/zrbJi4udBgj8UjkQQG/NxUpmTaXvZe9OYTDpT
uYhHkabPkHe+rMegdgd19SVSOrLo3rpjGIbtRGvmsuQOrAimiNyQvSkQLgmDs2jCOaJ0ElXbeuLf
E5eTilVMUhnVmoQAG/IWF1eBIe1LgYPqLIs1yl/I1IQpTPTm6HpEhNl8uZ22VOOwokYDZkknyALV
5HPONYxEl6rFs5kD20tY72Uy17gpJvMNC12tTNtodSNkfAA4uXNqTy0MP4wt904GgDjyGlbPrssw
YDFxd9n+XVNCXTMN+N5MEUa8o80IT0+dlKEqS2y77PjyBph+HuIDG/+XNYQrLTU6br8MdwP7oGui
35Y5NfLcCxM4UpA+SSRc7cBSBEL++lcyDlUZlsN2brALoK91NoknH4dmNFehPUAUDKUrpDCXCOBZ
4JTKMEiSlZL0Z9SXeOntb82am+gidt989EMTZ5d3H7AfQ6++T21JgK/SJJnTJLRu/dPGccifKu1n
dettmq0cSEZdz+k9cZofz1QaAKRtDeaq0Zbg8xtX/kUhYHSU5kw7d2wD97POUY3jW7mOMcr4bbWd
yPa6XYasZjIUvKj0+KrzVzBJn90xXPbbNsTx8QFtGBIAo9fDoiQ6xZIacXo3ehrmywn4N0jK4HYS
+aOMkBuv9bjkCY2+BWbzIELZ7Ix37EiGWUDmIEyec3nwn9nadxL50y4MSdvXWWdViiwEmQcJgxF8
T+qLQ8Wbg7F+vrKXjgtgZFZC0uGpma6I9sa5UCrbais000i1A1WvMjWHP9qXnnT7grmgV3i/SiB1
HPdmstY/N7VV/aYdFc0lihbMYtRfIHCeQWvtXgX73lX9/N4POiZccblBwfHU5ckqPRaHvLFEUc/c
eNdzrMDKlp0lURLQDwjhidlO3Ja0zgIqNmugQNPAAv2/f8B5lvQRq4/ICmFB6tOk52Rl0GX8kI4X
I3fPtPBcDuHyi8lacsvtBCOCoYb/2nQFP+ap3OsZgs1TrTEvLVc7u5ibLQk/w1op1BnE7tju84SI
4RZ/JFPx55rU/CVkDHz9UGpkoQsmRLJCvkOKNLzL2sWa5bC5pZ8qib/5Ej3WzPO65ilQ0Ji9VVVF
dq6m/P+SOhvIbXDWSeFVpfxvvA/AmANQi/Bma68BTl/os8Dn2noV9hu7b9kLvbCDURFg+FnthSkz
NqvaIdgrUozzWnKujqZv7MJO03aApuT6ZN1FiS091pY2PgL0bAcz7R3ZDiN8mNUUo68RF80IdVML
5WpI+ETplyrUjcm3Qti1Z/KPw+OfnUq/+QagQ1EuIHFWTbBeRfzvct/xAKtww4cw1JHosY616D8Q
EvfC/j9Ml0FiSDdumqraCxwwFsOCMSsjudFy/7dzgwkZ4FZ2l/J5UB17JSbgaJg0A+e+AoQ3BhQA
w1zFg2iEK45rJXQxCpqLNR2oV8Wj7762GlH02xyQHalqA5aT+jUJHk+LouVRUqPdc86QB9tPkZ+9
2YrEad+6x12kUdqtKThb3M1GMVHU/WtO7foy5noS8nyJ4w3ekoJFkhB+J5dW8Dc04Qz01J1HDQD3
lmxJy7jo11qDwNWDrbGwKYIe0DDACqo/iWXZHXzC97lmuHZkEV3kSXsBnSM1ykrd91hvtJvArSPB
tOkqB6FhEAf5BTNFxhkHM7ufFoUIfgB1uABuwvXMPChHXBlJs+vqKDtiDFkTt6KG2ONXY+h0EyaO
LIAPQ42k4KIdwLKozpkkNP+p11qQ0ntsHs9CeTYPnyhwoECoVc3hd+Tuq7OitCSQJpwdCc356Dwy
5AuJ3wC536fbSqw2uTyhoYyqQRk2XzhJammagz7v9u1ntCuidjZVoTO5n8Jwqjx5d0G1Ja94jb0K
fXyhAe2OyNFvRSAdQaoEW1EAWazg2Qx9coltw1scu1dCcVViaMUcytXYZUN3h46HVHPERpLXJuY+
+RjiPIISZOuau8hoQZeYTGjf8++O3f7zvzLOspgCGpfiZ44JUWoMmvLJw7vkmcL4oT+ukVsQTLf0
b+oJ8wkYaHniIPgtV607IQYL0QAJE61em2YhDFxOibH5ShuVKvEAQL4SUwtmX/bkg7xIznERfEcY
C410TYE5UAdmKdJNpIIQSSBIh2MiWJYoYX3oiBTFNKeEZCKkeOyX06k2X60k76itfiXZwdQCDOXs
8bIE5bJSdS9kY0gbwbin/rC+MpD21J+RBfB+Z9rCNLamYR7hWDwtn7hu1jy35CfSmcwKKN+SqCz+
KNgVbg6fjXxcG/uSx171sQrXL87Wd1YcrqILkejd9vtLJhiYTX3MDHTkLTIfyLaQN5BmWalJ9bQF
s3FhHHd3sRhWmr0PLSDlufehPfjbg3jNCk0XWLhKO84APuhTz4AIeuUkYV//2jaIteCqqxi31Rvw
qLpTgQI0x5gEyu//KGYmb4zrcxRwvSjfEZWdXnKBtcNFJ+0SGaPus2wko6BhXtpatmfjYs+s1Chp
EwboEmx44ujIYbWu/cyAht/MMJo5pAKNfrkTIXfYIUro8rCwESrUogqv7GovFXTmpKNo34HqIBaa
8n23QSRXk1DIa1aobzz89phjoTFiOv1dHpnaFivzaek9BTIe/LixA4I+WrG1vP940Hxi4vog/1Eo
EvxVMsyQb7XHaIYCjVklVtcJ+FBDIDf788dpcJOIunbyWH/S5/9WmRwXBp47G3PzMQwxYHKbJR0r
dfUVhj8PYewzXZn2WbXiP9xwwDR765mTFW6ypmcOqBAWO3n29fVNNiP3GHCJ+gKJqX3hFbCNn1DT
0473fUj+nbXlCXEClSiPsfw2ahdWtzLMJoX8FAMm3gXLImA10/nn85U1tUUaVIoJ5L+Fcw6LDYzv
8EpY40Gqb5/K24SdRk+OtU3Id/dgOqLH8ime4L/r36nShv6IhwQ6Y6EWOsBJmrRajZr+4lo23sCM
PQ38aQ5KGPwouv0mbtk9YqYHeZuLxVlais/4ngxJLZExPohzTJWAEHtAUFrE7Uif0ek0rqWVRc/X
bsjovDxh+H3MUbQXk5VJDRF5iQpC7w+oafApfcbg5MS5hvl0Phk4Fq313kmZTOWb1m0A/0q5fheB
CHBXmKS5o21cxVGjNMq2Xx1D0Kx4MuzMY5zHJ/Xo7Eh1SDrvcsTZo1u5QZ+72GExKF7bHVQldNUj
UW4EP1sp0Kzr8GOuJwsHcxWHn7LWG1kcyU0ZRiqIORF/NvnlH49886CszLuRrdikld90CmzByw6f
37BpdiufVHG7jTopTapTb3YQ8exY5tx8h/Wg/h+VALW3Q0ygBrpkUCv++ivYoZ97rec5qxsK2IAh
qa+tXVGO91giL8kbbsKqX94uFm7DON+4bg6f5zcMv5NLbIh8y9IkbHLcLr8PIy8eIBSULKxHHQS/
pZd9HK65FSeiyJ5/NFmCywFJ3jl7auvGzw4yQRpkITLIBl8/605QKaBGQ83cRZg184PbNy2ak2W/
lfQQluEhzF15ndOdJdB+a5rmsb9ob4DkT3QoHzZsLnN4WLw4tDkTdZKHVd2J7eFJInVgxKQYwdie
90l6DcNcIJzpMU2Ui/HI8rTFIIf7Eehg7wXuU1dchD1m2EU5V1SuUYpAgVqEwhk/LIPC26Ee29+2
ae0JFRMkL2Y+kdnQ5U7MeIaGAcd8hFa7zPkvTOv9bGhpdUWlPPe2r9YrGAFgMINwnQi/YKPzx6Sz
9rYm89LuMNKhNYNOLxeOPJMSiy7o1BdFvVAgh8mqdADooe828qkFKp5wUsTM+WqVJimJC74zOwls
HlM50F2Vhd0/0zr7oFVr0AvA4cuB/k3L8YWZu67M/ggAhrlL32mG81p/Zvpi+KApesevuiBp7BUJ
stoNgjHNzcWLruXytSuGaTX3SRx2ksJc2SLBuTgrHLrRM/lE80+3/xVEfVpyXTFdzCgXu4sfFt0r
3b0HYp6aK+fjdb3XRn9gOpbLFE7QP4DPOeCG1/iit9dCdYyhNPL3mTEVTWgg8xgkDOQ+P6HwhCiY
DCbeUyoFavWpXQBQVC4i2A5b/GYDyRiThIRYT2E8e+ddNFXTVafQXj/hbwRY+VLpXuoVDVdktEJx
EHXrC4rGTj85dVdjMdDQlSH+Pz4nHimghSzOTykmlPE3yCEuCjV8Ma7UKAlx+YAqjpEPELCxFFvO
Y9+hj4g8z64mXZtmprueA/ocT2mnAMJkTVe+wOXGg6gHoaQuNqc3YBVuEsax/wvYGp6/FIEvL1il
S2zGJqJP96Slv2jxTwq4kdqSdBPRVgLWMel7hwv8/Qf0RvFUigy5AXldieH+fzpcFDp8XfdzKnr1
1soaY7M9IDR7ltJ41ih+wMscjOdI90nKY9kIBHiOUSLbcl98+z0hByIIBrxiHnht2znWOSyA5rPP
1anNbmvGEOLKSQI7O548w+UUZvyfQ5CDNl9drfTjmZIpRC4zcS2muXwYbAP74DxWpiNGarj7FRcq
ShcVws7P2Q1CK8H/XqYej219goOGg1fyFBTYGykcsbK5ccNZbNSt02jCgEgqro5VWW3NgceSP7Jb
AGELuLzus4/P9No/5USBFXvvewoeCVaU/XvBl5ZPQ2H+ws70jrOo8Kt3MKI4813/Lc9S/yJR8qUI
b8ws64FrQlPWu/3yzFDYSZobRHjicLaH8ea1oaoJ8kkKJSwcwtM0I6HczJJ5ppwZXNSvcFJNWXrv
E4ej/EANDTl6vyWGyYdD5teAFMb0aBpsGi/8WYrNWSqigUzRyb5oWvuy15aZJjEKBjgweS061WsL
HAgF0EixSZizb0v56TjGoGLjRYpegNX+vrexVUgzI0j82XJ+2f+dDiRW/coUbdm74zW4P12ts/TU
9R7L2hW+IP989fig0CeMmcXNAZG9sSFZyYpweWW2Kjivn+66nt/UWe+HMOHc+30ofRskxRD5fzZb
tRuoSU8keUIBVxtEcSKyxx/YQ2v58MDBXSu2JuwkioTJ6ZWdU4wJt/bYGmLuHJaGG02GbchNYPT8
V8PiEFWbR6PgQC+dyt78bXL2sY3aJAr3ZPTqTCSAR1x96P6O1gXEpTxKgqYcTfmAe8NV+VDn86Eb
5+2wKf7g3Q7iypZcQEg/cHsLcs/qAEM1edEX1EBWlK529T+RzUB//LT/rI1SiYovIM7xSKhbocav
cu2k6mSvJB2WiSk8teOq1AtKKa59Cx8NubyZVQFV5eqSWflnroSzQQpiRP0GhwZp3Eaii1qf87Ez
m8bmGx25q2eZZQkD113IggaKXnFWAYqHVrdxa2/OPWJVaeI/GdjDnnHdISvEWBs7U9/ijDQn79cc
23LKdMzrRAFXA5n36Sn4vnn+Q6LdpZLhV3vS9eKpafnipayDn8O2DOt97CkUua7kCXBSedSrT5dY
r5jYlmND1cmGRGgSvqvwYYO/wTACLOMLHJu21V7+fj2Fxdaeq3gi02TBds1pV71PYiEZPb15jI/W
nJpQogwqEJOxa8VgnnajgWI4IvMc7VA/gF+XReQi26TJevwnvoX/5kICsgEaUReioSoRly9wzqZ0
52KCyyqoVddruWhDUb6Pa1VFJuQ//xuBdA0MOFkpZOvWn8eoHZ7X9v8Q3YhI/v3wnw6mLozd87xN
FBPb9AsyzSlx4E0ZJ37AaE95rwrupF9hSmTvHgOpBhjdBm4N/RevJsRABD3R//rGRfMPBdO8jdc3
jC8eJUK/yxhj7hgeV0LLnYoT5K5whH4/jZ3XAJIIeDyQT9ynYmhpGmApmmyQ6W5g5bZxPojFZB2y
sa8i/zqgPX0MlTl6oZ7r802A8RbR+bE+TymvVwtxsVppeY7kjN4v1N+e8qctSTEa57HMrxlGKzqE
/niFNLByIfKE4I73Ksua+0giWxLGNvUX4vGW6BrzsqO6lIo1ynaHLFUoXF/K2DVTOhsM2iHsq3Co
7OlmJ3kGM13OwS4e+D0/j/Z5p6vFOVR0r5oMceK6lBPb3zOgRkYKPg2ygzo6FG9FOktRiwNlA5UM
Fo8+frb2gVs7QzC5mrLILyv+JduB/9dRQ3GL6BE07YPAattmefAhtjS1nY/XdFgoO+mWK4Izgi0/
XZH6brIPB/RAw14OKKKccpGX2ET/mWvHy2JGmULaC8mC65yIuemGzUBjOuZUCicgQQsmq3RVU5zZ
jCE+dIhChq9uzBoV/nRaOzgQHBOb7gJ7TSnI3qi7aqkkvCt0Psq15/TlUHqYLbfMF96FFy0sEwdi
F82yWhmdHV5LLc/gAsJ8g18Km7Afyzt4XVd68CLnpiz1heczWjqOnnFSwJU+DOJl51NgvlabrOdj
U6J3cLuixfY4OVZ8y8JJzCA8ZOQVwgmC13nyUi4ZrF8z5Qpqa4pbz4Nmr6msELh4ArTAuiQ2gMHS
BJy8Bw6TAmphOfJhMq8cP2ACXmF2jQLVQhouTDqZv9x/gtJpY/NvQVAJ/9P5l7qijUwr67YuIGyw
sEuBZA1t26+RoS8MGyVIWPF3Sq5jRR/SdpCfPDutc3BHdA+P/ftc9OFU2+LB3+xTqAApqS6ACN9F
o02iuKYJ7uOsyeuRwdjYlMyUmZNPvUl7DOaWry/YVfwhH6mDds9PFiiKhQ9n1g7G3+7yKf4qHyXY
s5w8AUUu3uh3TyT+eKrxSyCuHSsqO2BmpVZJonq3I4r9uUnKHq5pTakVEg31lZTdNHXcTcROjxYL
TioMP2gO5C3fWQvPYq6xx7Hhfo7Z/QA6/a9ontSJsmQ47FKFGl3o6paA3m2cXYIT50el/aOf40Ha
2tZx71QVRJ7pG+hPYrWRIw4nojY7vdclUI2/i1Og4uMREMm/HfdQmKRH7aJizz0Dv6hUMLsdXSmJ
kv3WeN5TXtxp4cHwHRcnaB4UWwdcukRqndKvLFw9e56KC/KRlDxyOEJJuatY+cn2xZqZVADei1Zk
zMtAQARHOmTTzqF9yg27ifLFp/vfUvxKM9IfWNQdroBSliQodMAwz6OA0AAtsP7yjJDX/+QC+TRU
wux28xK0S+aLArFqt+c3gnnpIgEbnz8KXWuprUbD/CtAsP5UyAYRmEH0Rfs1iFf05fMc9KbW92F9
cI6n42fd5SnXREFuD0GflyCDmtt+CXJs9gWuhQA+myLxxLYoaPwaCtwKvnOzVgBvt4+qVay+BBBd
3kUd7HVClVGH/2JHHGEuuNZEExJm76SKfk1od3EVVQgin1Wv/oLdZ8J1cbkJpdE+9HTcCBMkHvca
fIJLJwHfHGAVtbtn36eEHZoQedTZDaDv8oSFYLiAAHCvrHM18gyqDqwaFaZmVqxC01CeFX+N3wg/
ZOkN+W/NtpL/Fp8AGFJhwy+GVe6ma2jiWHxF70A79hdUBDhNLWmKKesMP9lEvMTMH8zIpW9r19iW
8Y1BQCd2HF6zA6QQBs8anCgRS0vFlQvKrBT229f/Z6uKplCfrAKFGTjqoWV9EFYDnAlHqvD+F8Ez
ItsU1Xx5AQYS/WJ1AKADX7IMleb734oLETmipHoGXm+ZSmnIsoEsD568UROd2DExkbW7CRIAuZiE
KKE7m6lb/cGnlMfdkRBqqOuxO4DxHIrru5dky24Jt1FuJ3RcXJ/L/i4DgVQ0wI+UTjg4kOLFN7gO
GNnxCmpXlV+OKq/LzqSl+jZoCuhI2VSh5TXouvmDDz5Z9+FNPPUd+1g0LOaX0jWRAiNq3Dzo204U
oVD729LpNZc1KIlUpVm3KgGSMJSGjiRMMteLF7MNj1+3sX2n4VM+4m8FyJBZzm15eatyNDxXfiQ4
0HlJujoLBvw0fFbVWFSoa+4oX3MKPbC8L7FELuqB0pupDcnfZ4dOPq0T+5lrXzbE758ToumMqiNh
lltYDN3/Mx2ysW2EhoT5NnpXejTUCEd2/L9Hg2YyqGcsoNR6YmskD6T1Zsd1RUN2TP54QFtgymxy
uoqJGKaB6a1ZpcOU3+wnKSrDDMQG7Cf7Kx4+MBtEkzTZVt1cgUTZETntQdNhlV1ZkU725kBToE1h
aa8veOKNrsGZgcjfWSDCnmpqLSxzmLG0YmLoCtPwPwKbJe74qwH/g5z6KzM0JXC1MVttzAhYkfX4
PTG7CZDtH/tOUTiGayOniJmhrL9T5XYnXixJU8538nEhsqjJH12dXaLtA06XtiuFG17VPEjvgJwN
bp+lKhMBrAOrEoj57oH67iROUF+QPrUBm9bI9Hesvpz7LM/EjnIhEbi28IOvf8lQgLETk8ajCHcK
ShCm6h3Q+BAIRpwxI+fV604mjY9ZViF9Ac/u9J2ZgdpKV3Yv+nmQ//Gi2fv5RJoNoDXvRvs6Xm1j
DO4TqNMDc8FZT8kBVq2b24gyXwOgFQsRIyUpJztAZZRRzVGR5Y6uvQ6QNRFB4uESTTqF466u7EPn
v/MZPiPi1ZyCjQybgvPgUrpk3dtiKB8SgsDskArJvd2gL57XjpFX8nDN4Wa5eTVV90mwA0k/nbXD
1q8979tka6PO8A8kEjEoSLRoGEoxxDrUrvW2mQaKhhD8rugMNxmPGf2WEUwPv8kQW8SXhNyAguMK
VNiP79V5et6Yi6uUR5VReiflZu+J8LiJXNuTpz9uiv2HQwqbrZUG1mzOsPspj8LfpKKsiSqoGVax
YC3CIIyomTutE49eTs7jO5wNw617b9Wg/AintWH3jVeDZhxD3X2u0g0x2Tm9A968A6Ar3V/2LIKq
LppO+9AM+Z6+utAE0NqkyK/Hm3lcDDDG3X+yeo8HSyP6d4D2cHqXwwYb/mFe742qciYHttMlnrZV
5NldYNHpjLQcnHTglJrLJHgAEOpwf9LNlJVYrLivYszuHz5ytIUmH4g5q86O+MCU1sykByRA6IS/
AAWKGCJP7s/gQu8ulbT8LFubS4PTchmhSMQYe3JJEegCLYk55rTxXAYBfTlH/bg1HgJ+ioXFKi5Y
j7Qye2TJvcmPgC20S20uK2zHeAXWzyjyYCCQ/dvYSb1b2UrR3sI8FMHXyZrcyNyPv7KBOmrjhWZ1
RK77Vh1gvc27F8noXZyl2h+4WlwAMi1ql1dughaQqu1qA45fx9g3cU3I2xfc3yr8WF1N6/JKtyko
VUX+BgII2saTaU71GGxLVcYzZu6SzeNv7b/jO51MS0JXWV8LiW1nshxsWpqG03uFfcevJtd3Tece
S9lma+HPkWgFtGqxuxIJdkknHitwLKNFNwLmAqZEMAg8JXI6/LW6rBi6LyQzxThjE9tZidbm4Alr
Qkku+E8qZfxoMSpOkgY2dKiEkk54BLfSOGlXCEOc8GuU8o49emejdUh4dS64ohLXSTpstN5Zrwgf
FHTAe7HDo8TBwu6MI2J2F7KiFRrlvP3Q5aSUeLpqWcia9hlawwoIKoTt8D15pAHHlFKl/cqx+M10
6A8cV02cCqP6aTA9AAoynDlXjVaIZuDGrRi2V6yEyq5kMZG/E7x3Jo0J0tU2mnF3zLHje4w5RkhU
k2XvC07RMAc5qB/0GPGSmGY2VjdgY71arXbZHwDqnjj2nf+cliDwWSXNMHjpU0Y3wxNa+i1Bew/T
djVtF0u+hGle2KJmudqLW2R43l7/zKLrl7mmV5h2QuMU1FGYBMaDv0Qocqq9oq9+5vVHyXJ+dEXm
qwVg/VHbUi5lvJe7ozDxEe4xTfvXtPR0X5dQQ39bYmjQC5qrpM5WDTnQDoOyd+kjhkjtnO1wkAYm
uFcL3AIv/yDmITnMemB8U0kgZUgJfP/r8bXFihnTWIMYFl5fwOl5uMXoS/rrOo7Vvlt0rS1Cp5xd
k+EhGpz9DpDogzMEbHJt7j+HihzyIj3lBFmrgwB4NEqHZRHov1/a/t8R5L1z8nR8+1cLb1w6g9wf
8DXWAJBWg5yJ73zmkVdQybhS4eXbU6BlK74yedIfT/2WcYG7afyqrODeRUYVTa2O7jiGh8IGCHte
VsO2MPRGqQqy2+qDb6MmCbtjYl/Q4W3OvI9lpsg6dSg2CmsPWaTNgdgF7Z02nlYfVxSdtG8xBjK5
jPGSSIv5iPT6ztXxEN4d+XcHfn/Dh6gc2xtkZRMWbMb8m5GRUCDW2OKQsgRM6ON3R79sjRMI9lPu
I3PswzGO7hGlCYt0LLqOJ5Gw/RTBGdBjS808swXTswhe1knN8DmmOWd2ZTHMipCgc0aGfFLNqP7U
PQToJAbLU0muDCt57Y2cR9C/UVs1KXK4zPBA6Cr8Wj8tId08mAHEqmW8HKbgnipxfHTOh1ZBzXuy
HD69qHFxGYdkL3h1Zk2JG0Lp7N/n6aHQw3WwqoajaspPB3/RWnWsyyNRsTK/6GBq0kyYXULeVWL5
u3RPosGrROd4ahUtQm+EOOvI/XUvT75vKe7/WoJrUD/YGAE5i2MdYJLQYKA0pSbwXx1gvXJNnMC7
F5+Z5P3VVQrx88HCarPd6g2yPGg+HaCaGwm4ExRLdpeR5x49lF/cfHJccKmk4cSGzjHoJjvDcJUe
1xPDTeaqxsE1Oh7+E93sSa4SNvlM1wr0l/Bnu+4u1NjaUSbj1Xupg/cHAmP//zqNNJ5IB4q5KQnL
BqjcpnGyFE/ao/8Pdg+SFgmZAWcEA/xOskobqUYEWPGPryo1OVE+VAyKxKzXE+jzqodiO3Mvu5sF
r6f/Lb+xopm6i0NqD6locX7SRx/oKQhA0eqzh8tbOqqcEXczbd5fxgdr70OOAtFhtp5hTs1L5r6h
oer4n7fH7KzAYa9oBXprz0v8bavNajVOL8KmMcI6NKFe4zg3SsEfcir0AeHU8Jp3tN0IyTYHPEXi
nhQMRRoTHt5F+15fzigwLcPh2+JyfJ3oyp+uxtHZAhvNqYC1qceord3e/aNTcCJmbYSchgUPEqWT
8EqKRG8482JehnTqyxa9Si9KLwouaQdTTt2Zpwvp15O6Rav6P5Va0S1a46N72Qob0B0HpKT2iNOQ
l7x+J2S7or0UywBTUXfwYtyvCWf/oL3PANLXjDMW3zCu3U1FlAouIUdpQKjQk6Ut9AnYG0N5VvNU
cZNOvl6brORWDCw6l0CvRyzkVvx8in3TnhZPmENjv+DtwzBoRy5B7RpvNr8B9RpZNtvb+aiSqgbu
Uns5waqzyY50reX0y5GOwOrMPbvL+RT1owE9MJwbVj0zV6DjRh9gP7ejW4UwMiGufT9Is1xthLmQ
V/1YMxmNM35Y+B9x8x6JC4pNRc5LMzxfVjtV9WU2URgoAbnEluZlTzajHyUqr8Y1WBSIEB9xqTmA
wBUYAn14FBzVqd78pE7S31OAYgcGG5gYkVhI4mXmODqH/oFtKq6ezoHM2c5YDRzd6QclPGwWoQwz
3u8ZWAkRNst5iY+jFYOWgZG9ZL6pclD75yKoKQNUFASqJ/hmB+keD1Eu+gPwfSvhtB1hKK6n+5Hx
hJb0ht46TiNuirh4tvroUqWhKuXuRyTS4o4HbW5GqUGGgiNEPe08EhF2XjlY00NYvdk/FU5bLeS3
6jbqDRMMjeM3ZTuPmVBYoGsJBTRNIEWhV76wN+uHB/zrc1RrTz7VYO06CFvog5gAI9Vw+RXUaviy
lvcJKTrEcIcKyRoXLHk0tZSAulew7ZRKrufugM6Vo5NDJ1LZXe4x6M6S7H5OaNyTEgRIPoGseisI
ANTzkAPmNiPPDg1ZH8Xb0vylomI3LEMkJMSGc45lBaqafrCwiG5urMUGK0yWh9KE57lAfkH9OlQM
CxJKklEgaUUWgaLwzgdTJhm2EX/xuAiInrsX+3Gxottx4G88BKGdbhK6HUSws4zIJQOsGcICxWn9
ad/0Bt6g6OF3R2E5uDIx1lR/3cYgzhf2o6mqFwHkwR8A8AIJ4i0S/v1ogir1shu8qjDrywJp68qp
nOEhItcyD9BXEnsJnwr8O8IGCtxh9D8x+hEM3gLk+y/qes45jK7Oi775TeTZ5OiF1TkWGfjTutrI
C20NivP/93TH0UIj5LSgRPQphZ4L8v8NnaBpGaJ6JRGj64AEM2LE5xD4WLJ2JZveODBLz0jcopYR
NPJN7qrOH4umPhXknPeOTgJiyvtUZIzKy7yqTW7R+kjXJTpRNulq4Yg5G10PAh7rSypUwQ+smbAz
W4kt81KKzcCtmwiAMyZVaJUoYhY52/S01NvzDYHG969/gpWUN/3S4mnpjeqH8IYUF1MfN0bKc6sp
OfVlZ5BfEIOwJJMBEosdiDZDSVcr+0Zs73CQMN+twVFMQ/1ZtGswZUgjQ2V8v2CWOFcgGvOlCV1A
R9hc6UHqNUoxumej3FL70RNlyNCN7VKXQRxy4UGWAG0sAeep3jFmlANNIAPBVwQYllHNGDdhqcIz
TQpDpfpd2jD4XxojZ4LS94XlRpseWulDAsos3Iki55d2SEruu3MbqIt9tJOrHDbRSkogXtVWsb0P
TfzwfduTo8VUmcNQ652eMVHuh/FXRRSwklrkEc6CrrZjUviSBZAhrSKonm0yzOwrawe3IR0508OA
IRW3a6Ka58iN3euypfh5Rl60sECK47WoltKSEesNyUcd4WNVbjlo/S6kuwWxumonG/lhsMZaVlLt
eNSDDLVsGHBYjzelSyommnvGchrhLoANHtM7WLY/2Tm6QibjiqbvrCRCLQQOt/TpfVWpAfLz+95I
0TEaU7KrTy7gMDZR9dMDD09YnebjecVOx7RwEApcllAEd0rc+yJwPzf/WtVTrJtUBA/AydKcBUKZ
FZDgMimlP6oqJehqfq+ft8jTh/jF+F39jejzFZe1zx1poXngDEXsR0jWXzY0wKlohZ7iijC6ggQg
WvD286oBUhEreDiy7VE/39SkYKWeZjXn2/6NV+/Js3AZJUL4ERz9JNHLIdEDKvv5dyje0XX7+DbO
6R9I2A0YtBIyk5srbUc4Z3TnsZ/rMvMqE+saik/5aYr7G1TFiE1DwjbPqc9qy0k46RfIDt1pb81L
CIHMHOQEJnOVTf1XHVF1yxo8gW4WgzILX8NllefkClT/YhXaNowPLQtl4MKL7dxx5armPWY/xFRa
hELBPZepYHzOldtS8xZ+U8uznbAiSrqCS5hR4CIYpbtUB1056trMeHKlwNWr1HxgsYh5o16e9KVS
uAasI2k1TnZA+6PMVxm9OXClG1rcrmU/JVul51RriCPEr7NWf9MHAOG8gUai/OqFcSt585vWDj84
ADF8Xa1ItV8ii33y1q3OtEhjB/wMuNHwZrKS0LWVm3GjqS6k7h81l7Kya8wyotAcqSayq8KTwbgu
cpezj0rTNQ8OiTkEGDJISUPbtA+AAstUN+n1DSn5clloQ4mTPiGS6RtZp1t/zTandor5slzQbZ4D
8e94eQbWEMH8se4UGT3BgNubZax/xXUx0tCT51HuI/s5pmhlqnS1FqOIHHz4QZl3OrHf3dHFbyNC
iliQlJ2q2ndUToKssz59Vl6tkCn3IWtfQsiCLopSqnqAumurEaUW+qgNxr9FViwdgdH9+BhiRML/
pM3cn/jQTrpjBBMPKc8ZK/kDuMQGUg53+f4Zmlk7DR0JhxiXHpT0c+hurqkgA3BKmCJ//cNJuNPr
qSxHLJ3JvlXDlU0g4lJ9kXczfxuo8J3PKMhdO94sM9Sc3JC95GxpXKcTbm5q9TidJyCNW4gwV/6a
VDaVwGhAgFn6u3piXIYT6uu5k7mrmDW7S+TKpBkGwk9Imz3wRXrqR9H4PNAMUtmNLzR3fg3UwPX3
SfF0TSV9XXSSKCo2yFHQZJTqYP/swU05K/ECTb3udgh3wVt/pylfAHCmcbmtANxANdhLBIdUt7Tr
7SJcO3Ca/WuD3ZwzGgtQUrLi8jA/U721ktvxFxwvl77x5hCtIV43feX7J0aB55sRCaZRJ/rDhOAo
mnMIs0B9BXkqnEAQZP1wtNGl/L6UmYzl8VZ6ccMeYHgKMDwmmCu8cRGuvDPz57toQ9ved0gL8a7z
f29reUXV9Gcm0AYf4vDv5JrAxOopTSp/i+XgMEWOcBQ0Z4HfPby3mKsnY8zOaGInxGhF6psr6cVI
7ULL+JZUItxJTTS2x9obCJWHK+b4jhMKY6NBw1E5OWkYRf4AThA+BjIv7A1pM+EIaAdg2i24pI2e
nRQedIwxLtlOtEzu7nTCzGqCJKQj6DIW/2QaMmNxWCxNKtgL7KlAdAt4KsS72MJIU18AJqufuinx
kjnh1BQeDgyrnZITzkVVzHoQlyY3aXdG3qR8EywVhvDY9Zjf1VHucxtk6+e/2IAA1aOyR9EedIT3
jbqsSccmVsE4kKMjSjoVSvKcmEEm3uX4iSN1YrgWQ9hNRD2fyHSc/s8/FiIaYES/mZrS56Fpyecb
HAcH5C2FZF7wE24rGfMp6D94b8YLh7fMudlbWTbxnTxtz6PBYhYYk4nrSs0r+YV9kjgO5YHCDhrZ
tcv4zBkXPTKOsIbleJ3kLPTYCv/CXmvKMpt0uwEQQHL3q8EsCI5iUjlsI8mj0cmoYDjf8qpVdV8T
KYz8GPIolBAJfODxmQDSlvJWZDuaJemcDdjG5D0FAhY7cO2lDtaZmWebxm7FScU+P/ujN3zpcxOK
2G+FBtN7otbg6MTsAgpFpEIqHnHIT6lYl7nCs6U5Auvyy+xihJuFpqjQQnKILqMkz8ZEGRPb/Tj2
/nt+9GvTjLWYGpBIDNi6ZK4UmkEiCzMiM6xxctKWJrNdSS1bT2zkqXUF6+rW3z1GOHKdRwokgkax
Fd0dSxYQKS594Fil8s7X3JX0f9/tuki17PxLjR+MXI0amW5Lnha86m+O+DOPICqZ5wTBl+Jj3dHy
iG4GaGJMWidJCCjGN2ILeLH6i6JnMa1dPB85twkNRt+je63cHDbHUymfVU0gkQaQ+04tkf0B5fAP
uF6LnrsvWHFpkJ9rXnsd1QzVdf1M5BpDYutTb/7BMC5FGFFo4U+Uq/BLZWZwBEARIkHiTnMERB+V
DEhgi8UsHyevu6mqLWLtPtysKB24d5tcPu/23vknd5L4mJtB12V6UoR8AH8y152/rbN1xLBjajII
FlbOxN8wQzczx2OMhj5GmNCR+4pbe6v/FaYCdhjwHjdgwaQtCO7X6nsApKyv5XMjhM/DG65dgebp
jwsAbZTxexfnJqbF5vi1PkYb5Th581veYNZhF+gEGsYquSYtALpltgtF8KpKh+3duWKACpFo955X
kuNRlVqMH1PCfB/rjkyNjYKFOa3Xq291qhQlvx4S/yw0mon7ZppE1XLYwBzEM3JxZBRodDyi9xoJ
gC0ytv7xYBDKQUFGbz07iaXciIv1csZQBMI6u9eyKEJl5jdprfnmFUypD8AUQ7taEGroweA/oP71
cBBVw7BmPoesXGR+L81Cgq6SkTAxArQI4wOjMkYex3Xf/ANzgPADKdCLPx2ZiVDfFdmHoqr95kaW
K4YzYdBxcKuEfBi7fCaIOBhKYFGwnLLzKW9/bxue4WjS53QTr6zjZvGqRXfR40TzNdwa3Xl359lj
hAYNr55plDlrWEyTRBnkqGZP0ZnVAutc7YBkgZAPs/gwmyZBwbJZTPf4oJsLSAr9Jvu0e/3LS3Nl
6EJ6N5uPskM5I+9NOaTpMD1ly5icDUxrdonNX9RwfD7k3No1LJeYgNUN1NVLpC16azMZomeFoclt
REAC+ckU6kNpGJU9MdPNyCGqw5FSSQOXnUHqpOMWKJEsWYfGjIHBtooadJUTuY+TKWtLeIX5AdFy
6WbyyTkfhGyl4EqXzxd8EogWeyC7i25RYVU+lmt7m0Fz/9E32nZwwiIeHKrNZoVTa5NhA6GlpfgB
6WNwH51bErmyo4skPJzjPwmVBFSj54XRQn9XPudGT4ej5/ZTzAJsAWUFhPOCKGPtTlivxcZupbOU
tu4oZPG3T/4QMWyfDgdr5iktndnVtMC0fSmGE6FCn4vYgZE8g+iXXA94PI+o4arXqgAsvYTTu21+
qlCxUnWgJ5wf9Ad88w3FMnlQhM+7EuKw3/SrRegl9lVkdIvRcePtQKAY2hI07yIL/B6jDQS3aSRi
X3hrYQDE+M+Tvz4+aGHoMxdwRvRvZCHgLQdvf9EbzYFoOaC8Dq50PrrLNK4q3gXlSAkOYSMr8MEE
HrqBZcVZz6k3inTIYTJwIB0jJG6vAjSNzvWhvcBgWBxpf0qeWA0da+pTJXE43+DMBEPrIAM2vcWc
BOCyeWIlxqW9GDxp5u7KHCfMiiTirJ5thPUFm+8g/Ne8bS1KtXmsHky6Fbf7qqsZWr5tuViMgIU3
83X/dmfvayCZrySjbNU0coNveS12DXCfl1Kh4F1dpP6Y/xPBukvExV/pUHssQvlTaJgVG4fcv69d
kWYIoovHmvox3jldsxZKYmDceVnTh+dZjgep0y6CvzjMFdpsQPxPEXXYbEiLwWWhxQHB10x5Is+P
/Awiwsa/z4m86/hjmknnfhxkM1aV5stwc0PmN0qHQUm13QZLZ4FdY64ytkW7yrdFivTSh5qRQs68
W7imyfl4qsG0sf9m5azLrz8fjbs1/EzvYlglRBfTziqT+OVs4S+opEzZ8v9TOwF9AFQPWqlkl6qL
0UTIUlOuDh19EU0tvQlLwlDJBt97nGL8CyRKRAn4UCWkBjWZAzGrUH+sJ1nihcTWY/y/em/S5B8A
O0+hv9SP0BddeeaHeQDJhwWCYd7lg/SQYw+YaaUCvZlJLTBgvBZBwAIheDKSVRfD+rrwFrb19Xj5
/scy5cRKKoo0rcVj+NIQY0o9qAXCP5D5iPnXCg5LJSWjyd1JFOD7jXORZA3hH5c5Hq9AMH2i6ntR
cV+H2hSrGMQ2/ncIFbxv3v7sKiH5LGRZm8DRTluiyAsj1r0KQwkgq4ycb8lXyYrnjR3EVubXuQ3h
MHdeSst1HIu2NIuTdN28DXCO4BNZbKwZ1TuFTJzLmUkivcuE6kvIbJOvbivF04XtyBTKsnxdlC7G
83SvqWM660BCOMiHfrzmeu51+c7mQZ3GuQNIB4y/J78kYfQpPwDumCq81aMUJtrlF/ZfRwmml7mS
wpsx8eiMsRcSBhrHzCGUQy7SUjJcyEb+6gXSN87kJsqLVo0bg/kZ1pIowoLAqzaahE13P8zT1C/n
ofRgmTGB0Vi0RlgU4KhM4uwWOEZRCIJRTrQ/+Dix63w9/Uwcnk9eQfkKX69mJ8Ir4Hbua3XagwRF
YW8eRAzt1hUmMwHyzfpU6FOemZ8ChD6h7rGdYIxnfLfcdSKWvz9nYusoRUQjhDX7CldTs8FVwAg1
BM7NUabbYa4PUXHlDhOXA9mLqy+US1xKVi84xCdG7c4nacZMTQZtlowehBnfh2ICq5+CZKP4xTPK
Z79cLKYL9VWzidKksNtdMEUkkfu6Liwj++/zlRGvfjPcN87lTQkIPzpUbMSZ3whf7iaAREXKWGUo
QLy8teIxThTkTuBNFK01tkU81tjKQ+YymrglV+WCY8536bYozYrv9Kxaa3Grpul7PWiBOl8qeeQD
84SnpL8diJU3YKQEQ4LeiPBevgFKik5oXsAEISCtXYJ1mX92VNBk6jR6L6B+3Vlo8oiSOCH1EX8R
/C2sdDh9IW8V73wKQ4JD2y08KGfshuwGT7b3vFv/+841fkkq4bmnOarZr3kZM9rDWEAAuC/eFqNC
KHQVHC/irYqjYXWjoW/lX07ZnMls9JitfaE44UKu/37N/KUWxgS37KGSyj0xLZmUgO5/Ndd5pByN
hUczKYV7sjBFIO9F8F/4ppCBlIihS1mCOPlwARO1c1E5j22p2JYgz/TqK/JLUxxOq4MuFnlJ5yt2
uxwl7rbeaSkNw0sjNn3R55d6/UvunxsAZo5od9leJpwp3oOy3kPyHJ4gn7Tmg82WClH7VUOn426W
AjWrFyp7zXyctKtLzrj9KElD35AlgytKgF8/OyNMnlpC24UoBgE/wsF/4bUV5JOnFqF8iFlO+7HH
fItEsDC9pyqluEit83Y7/uOS4JplPQiPqK5bJZgvbGvnKgRBiUg56ownySM8/WMXpMZ4rZaWsjzU
c0f2remyNC8cx4uaTHM05zUQL0LDKcdync6eSjuZEp5ya55MB0jHn0XocanuHrDO4/FqQNVgWzbE
maeBDbs76GFce0u76YuAmsfAezgLsb9F6FieInTqvbERFeBsG205a/aOdy6n9uBy2vpD/YYapVsR
CI0gzvDNAhJlXX96ZWeVnK9ocdrpouynp01wEqbGPNIKZd4IcWUYBMNr8wvR5sQiIGx0dHmG2wSb
wdcSFKyPUBLGihf0cejhD5LGeW90Tkctbu1OLaIFJVeuazAg38LU7cggK5PdaTWAx8am4fL/WeTZ
L1wxdgMeIbO3sco+nt4SM99a0zQIpaNZc78YxqCqiYMROPCKRPuGdyEgO9ZrsOgnmhs58j+L6z/5
wVnskv39EmAQRF3DBPnN5I2439Q+XuP4pww8EzC7+UUgJY7yLrFzUynHTSGoSiPVPhn/ytJ7t0jc
vt92OsYPjGXjUHjj5Ihe/gr6P0euSsvEed5p9k8oNKyOvj5bc6aIvFL8KQ9J+YANRUcyn2MA9kme
xEf5IP2SZoRsmj2c+IckLVCWGZ3DJlxWtBT5nhHfnbueIwS5J13Jnkbz6o13rf/IbH5lj8zWoRgl
ulD/vQLt6PSbEh4cN6Q24eOWL9FlN/IhezJp2ZWQhquhicAN1z20BUkNRdV1a8cjQmhQS6JAMwnl
tbNElk/6zGnCgz+IOjIUiURBDusN91fP5m9kLTcz2mo/5wi4VRFSqyNHyYv7nselpHYSnEIU1ITI
Njyg3fRKVBUz7mjxMreG9+sEHROJED4IOz24vxofxbthUBTPDseVSljfwgOB2ZH7gpO/NdyF47us
ql1/Ylem/hXdvUiwrq5PU+/j82AxKUvgIwRqaVLSALEMrwNU59hVLy5eHYLuZw89QzYzT6wUkGTT
oouhiRCaUBPr3tqouSlUodps6kr/gySG0KmgfwSegndxeWqtM9Ft0s15PvIt6hi4ncI0lf8oihkv
o+QYAqlxke8FhluInzzjCloxc6xiSgHktYQ2SV5+8KTe24U5o5qBGxKHaogpVbhVBp6GUa7AFCNF
yxnmau6kIUjnpgUUumtGtFW5bYRJzZPgWtHrm9Hessx0xRJaa1bHavDSkvJkNnEIpCe2JblLHkb9
9LSZQTehIXTYGYZgAwuWrpjQPpNC6Akf+3SbZNVF6ltW1YrVOp+fY5gVp7o0XbXrxhW8pvhFvVg1
6XqWuVejN1UwzOx7w7FInlweQ0n+yHjMdZI7KpxgbmfqW3lkEHoNg5z+YhffYOC22Cten0u4W7/9
zRl0/Tz69pxQyNmuQFQuTZ0VLeQciJPa50yo6FS7+IaLuRdHd//+9Sdf19IHpaDrmVrLR/97pwh4
J0/BDamgkiSv2cG/v5QaR8Mt+L7h42QewdRVCZAkok/vo6oVF+7mTa7z8EP/AnUSScIQMQjD+jE5
auomDrxFI09t1Ob5yxxiLiImLwPEq/JkBHz7DSzFS4GKj3i4LFeBaAQ/YHDO6N64AVaKiveMfHls
ZtuoUDXswQgVnaeZeIj6N4hKGeQ1atShFlSJ6j91MS8VuWFImbGUJXAd3u6E362qI3D+tG1CDAov
wVk9NUfs0Xh8uMcG6VxTF6FvFtLh4hbD6p4JZWLseDmhSMbqkGV4kizkOwEg3auVKHWhC/iXAo2f
6Ha6Ob+RhJ9c5JB7QXN1lu/VewYkBmCF/wO+VVlRiwvAx3IUACJ9wgXQzs6cRkWV2sSUSDsQkLKM
uvwwHGHSrf5XLTmpqmrB6hrOl3csjuyuw7G+mPZGW6MMzwIWw1IP4VVMGXhLkV2zhk0FNO8Azbzt
UKb3JHAMikU2VUZZQDLi72Piv8IrrWWD5IJr19fQuyBcvIzsJ+qW194WARg5Cyd1X2BeQM+lR4ol
ggO3/9FvxGBLUDOGSkhhutQgyCg/G/9WKG2hvLbpTYpYvQY8toKyL+yVq+N2ASeb/D1xkZi2fbbS
xwyNlqdZ6dI+Dlw2WgBe5wTgaLFo3Pw/NaxyX+VGyf02J+M9Rh1jnJ5q2BACzJuOepwKrE0SpeO7
/XHDdBdBX7ES4oYF1jQ2sIchbRBRMvyHd/E7md7vGSsW+xitP+Y8RTPKUjgtxPMdbH96xPQAgCCJ
v22jFqGNfKCVVhcrz6czywidAqpQXgEKBKj+PtkViq0UlpSf6P8T13IfsYwbfNwMGKnZ9VZpU7fH
SFx70MI8Q1drSNBVNgGcYOtqv7iNCojr/yZn3tbfOW0HYLRGbpvcWauTnClvNUYGbUWXlcEyPwOp
SvQ8jPIzOXOkvu7rDRfRF/B7yzLFJ98oUpHAHb94hx/3H70HzvUyYywH49lZUFoC6F+mmSwOJxH2
GvxWyUw/cuk3VrJ8Df7vbXX3awy3izOQIUNcVe+OFoQGwP8XW3n97221W7Z6ZhfsWOzTL5aZRSUx
WWX8AY5l9yOBmVP6mK0pf0VdhpVc45nK9nV5AkfUZT2wBszTU3+kTXvbYxozasmH7CKC++GKiVSX
kMIjjaomB9NHbClIjwqv91ojF6H99j+d93KOIM9Kaja0ak83OQmJCeey8Wg4OjY2U4ZIe3Wl18JJ
GGG9mN4v0ZpKpq/doRHWoXKuQFrxA4v+MvkiBEcFMrxW9RdzV53iSieBhYXDMGrjz6+0CFVjrQHY
HH2/UGvCotSkao+U7pRV1GEbhyjG9Zt+HW86LA/u0dWILm2kc7dmkrPH43g8aqxmCEcP6NLz6Z60
aYh/dToNLWBJ8zFSfZ1YuHtdL7QOavzXopUiNkL1Nzzq4i9E0+3S8vRguhfv5VkwJts1DvnfbxVe
B1KZrThvc05BTq6D0k190fBU1E6j/V1++Y6QUKk+Sq1K8sX8FTUufAtDzAOFQzj2tCa0WLL9yXa5
yUDpE06KjryAaLtFHV5ES/yn5SE/lx9catCCOFJPaw6vLILGJCn6r5kJy6q5fkJnEwXvFz/XQjyn
MYPqEWRJBveGhvzJI1BsVUHdIOZOBKl7TiW09zOKuJ1QgykuX+gaal8kG/3HyMfgnEVqzAc10TLn
Xx6TzRoCmYfcCLPLg6x/3Y6sgvq8n4zgNScF3RXE5nz/wg4d2Osirj/CSP/HoqqS75RO3N4lRPBw
ZIajBQMakBw3g7wgkcELZrpA8QXA7M+JILT3ORLTdVUfMHkpHbE07NLZk2k7DMmuchP5PCt8wLhe
5tcT2uy3wInE87Dmx5Mvur6J1WjDC5uK1yp0OGNs/m5RbYujht9sT0O7sbFVzY7CxLdh6m+HtZBL
h8a3wlIKbZNCKzShHFah42ppSYi5dd/ON4XylfulfwskZGlCGbpUdXgkabezVM+9NsYcrH6MRQJW
rzs794C5ni6h6Vtr5rpzIaXdTpkNVCrGaNENekPp1wYhvg6aKLMhaQjepOw4mH1tnBKnWGJe+7z6
jnGpggV4UnAxIpfwMW9KWJZIWZNBkJjE+rFgcaLL+fXUAZdpy8cczOOZ2h7N+rjrXYDvhF/qARDY
txuOv8t8/mnw5T4v8ZGwp+tKVxaz0qPJfsutO/mf7g4EHkdBLCjS7vg5sTFCaeKRYRqjPbXQnWOU
Ke5x8a5GVP+5zLud7rS/Z7NBZyD4YqM1YsQMyYqYOjcy13v9hA4K8jGb23EjkEYez46sbMjftYDs
uTcwnTZFU6WpjOUg3zFSpMdk6Y2n2osvQE8QH+dwcbL97rwVhe+Bx5lM+JzLBTNNmwykK0IVVx66
Zf2eBDXjGJmlwH7qjvdLCtCwsYchZ4IZaMZT7OeHZHLb1Lzw2qB206Ndl+AXL+Oa6u7CR6dYYdgQ
x5jgWiWIiFYCHZ8rw6nqq4TXBsMoY6qCIWoQnRFaKDub3co1LJxeje+MFpkwDIVn84RGL7ft6dh6
BLZmF5ycRr4ZhYLSaVEVXebswU5YMRDhdvg1TapY23nlMCifxOtofAXsNBD/4SU28Gncqtq6UtKq
Ge8Ck5LICb1CTob5DhE6IRD0s5jHfH4nGkGwywYVrYD43QV9pHAAG7H2v/PD4/7I14R61Cisjvvn
V84Fd+pqr+pAQfhw5Af5doNyQO+RAvS66389ZgsSA1wBq68qLQSvOzk5AT59T5B8DmNr9+rQk+7z
wh1bwQAjQmUZ/m8HWAbxWeUeabeCPNA0bDT0POlG3yl/xMSlL4RjFGqqabpmTG5dGcaMCcqbnkw3
7ac3uVSukHwKyBAx92QmXcOLVqCbJf0X/y7/8zNsc/6OFziRMwcttUJ33xc3LXjAZA3KYJHDg/6f
Cl75MMxEjLdPZfjokawOqLqKOpNGz2yiudXaww09UKHTsTrsRufyjh9KDPa57W+jnaodb8JL1Zdo
4/4ALcxVDPk2QRSH46aH4bN9d08niChUmc1Zi762fQ1086FWXY3h1KrCBozdsGmVMHN7JjFItBui
o/8eWFJgSCMGIgLgoTvVhfpn/xWOzY9Yld+SgiLHMgYw9khnTpiSqwRcKS6zxbIjZ7WcZ7kJoEGr
5P1HiaVvhj/fGrHRuVKsvGjwe6txca4egZs5h+8OfA0jO2xd2pP8bYAMOs/tHn8M2P30SKAcst4k
jP1uIL3uRtn9YNLY0dbU/XCjNYxOP00RaH/AHKsoFm5NWzl+m1HDwrN7J2Gof09neVDERYRpzunA
zQF4qrgZpM/lzE2XltIbSBjDT4LHnuXag3iQb2snWkQtnJ1v4yvU6r5tLgaV//ejUoYMZEv2MTj/
iNd9N2peMk8eTMc772QAyxvOnWaNlw5+wwKx9aJIniknClvqc8J0DvIednK/RKfa28o9shOBuBMx
HoAXNos6wuLPdQrmLBiKcuaaS5OmKBEPlv4CO+sRHZFXYxPQSPdwVDmuBWQlTfT7JYGpkxsXLBNZ
PIS1MXS6r66bjTXEatySaSI8KoW9NCk542/05MWZcNB36M4yRYGO6igo6+993m5TdTEVTcl7fbse
BwpR89r0Fbo75dh9+UicLXyYGgqG22gHx6yUutV38qzeTiN5E5d8+8jNnakgImVGU05jx88RKm35
TQfb8GxMRshEzhanXcTeHvOKimOo6gNwHH/gXJvI96xd3LuczLJSlZwPeTeRxQpHglWOZKpGuxFN
nNHDklKU0hf5+qkexyY4Yrh4trMpZJ6tm2wDHQ/ldXCYFJ5kWV89YNZSfHI+QFfEV03QoR3Mm4v6
af8K/2wZ4A4z93LhvWQgyNPwXSIzoxCH0657C/ZBjWtHN5JDS+eiIMmQC473dUnVU8Xqz8DSr+/q
62US2K7BfTIKbftJNbqAYxmO4cOgC7Isl9dO3cWFPV473KPRp3e3FUsVjM4U3HGwXyAA/tgfs596
VGHshpXQSEUYzVh6g5w35ZH2i5562TP75oToi25NLM94q4lsTBz+D9hTkjOOIlZIcNz9gzjBW775
nMd2cuswHwBGlUOU3SUIsKzQg4bZe3Kw3cgUBh/2Ux2Q/W3gTO8uIpaE56YMqx9GjY4wlioyT3NU
4Bc2xLCfBxosJsxFEn18bi8Z+gp7yyruj/7kZkARaDWnOBQqScvqBKzRPzM/yxKc1R7mcR7Rroev
RzSxZuxq3Bujmjcn+vHqjqgV1TIKjV7AuSTCXU8rFuMmt2+GAPU4/YPDk66Apz9PBDb8RalUd/K/
Z0Yjv1KnxSVWmZhsdgAMm7N1sjC6DdL7r0ZP/VhDrH/CEIYZV0fq21+D6sRktqHzNNVrI1cLFXpx
UaGnkaVqjiop6P0pTl7a2joWYFn+O2H89bnRudl76nlmvQELxuUUJqOho2hcU6W6wPPy/acTrfpB
tG8Z8/IvzW4xtHo9wFpY9vk6tqz8rkE9gFOZUA0M5WwvkXv7xDpDRTpI+0fYhHpb2tglJboQJ3nz
mgzGKCcoW2JvtBtSsL5bpBGw2RpGZxCxWy/0AlqDy/5LBgR0tYt+0vlqbt+E9UhL3ljoKsXC7f1d
5kk+LE+fbnkfVwUhKizjoD6JlrIDASsUNrl3H+0Vr96WouyMgSlsSER8WnPbYoSwxsqgYPLLOFdJ
0z+1//utouETvkC6XFQq1bEYSvfmoxsuVYtU3/NkoXY/mn/r7TP1rhC7P2Foe/tTnrLo8xWFSbpZ
ljjFZZCDbyF1y42yS4GTj+Zdob5sHzH6qdQeYmlXdWtAE1ii2o/E6PRSgoh5QVcFuf9i440pRKP+
pyUkbYgc6xDowcJfSSwzsZvNcYFUUBhUXgvyuwBrpXAt/+yt8I/k6iUwhWcaokRSypZc9LuL5fiM
fXPKH08bQurNyOaGnKV7FJNjf2En270Sky9vcEjBS0Ro7xOhKG/VTIEcCqm0myixyE/kTY1pR/Ls
jZBYbMXd5Yc+KvkzM2vg0oTDd+jO5HzF78eLT0MzjWYC4enPZgeA8XImZQ4qRY9l5PWy1uhwYZ5n
VuxHryct0u0SiKrgu35d7efiQQWdmGjjKrvPQOcb/hKQXCpr9g8VnZvh8D8+jLKO6OGPkCDPBJR0
s/yRDGQv/auMuElDV4zirbufCMYQeKZ5KMU92ylkhdE0w/CrlhuRBMvpqMEXv+A7hSzEWpBQHLjA
n+tXGSTf8Uyz2AY4s7j51k9STXKvwJJPenL2slREDAZnD2YytfgVW/xgMwokiqr273Met8XvmbXk
bzSwcDpWOvxeqtRMu6d3tf0lgKLnVe4FyyoQ6tk5kv3qYrQZVoy571nnq9g69/8gWEswySNQOKgA
1kn6/hEUcwu0DleKugSAMScyInyCwIyFh32gYKOs+UeHtKCgMEKL6ubEi0VH27fNgDWSpBev8n2j
M1ObnY/h6HdnHREgpFt3Rj3sRbG7L7+/5Wl2+mS4HVBB4IZgbo4xoBujKLNq5n9XKEfIRMyz6X3W
zEPz9bFoI4L8vvvzAOGfpJbUqpF5oih/7kRB6Jc14hq79YJQqLCcT1l8aIsnSR246J+mCx2MD87g
SUlrG2/PJ2ewLi2ra3F0wdsd5MMgPb+L9CLa9WbMluEAFyuzcH3kOEm6UDsnMbvUDyZ8ZceqZqr2
SOKZ33GgE6vCMLMpC1U1BzRpMrfaZZWTCuiAlxlkXe4gabZ57x73EbKDdqxU2pJyEzfuzpdORWXg
E07bXgdd2ShKdTYygv4bh7z9RuLcnGeN787tGK+HwtTLk26KVbV/n1mzC8FTzlSYRVkFIYGLuq9m
vywEMcb1iQOGAjOc6dir49Vjm48PsJ0VGYW6SL8BPbQVsZxPCvf5bv14pFHLTLSfx8j95PcrQzD/
ZFTu/KDXQQrFlsHpnlURsPacXOml+iYUtSRUYdGebcUD1oPvSaNSWkNcTcHvv8FC8JJdijf8luo+
kPfphQ70WkeijFmcGAJ/68p0rP0Y47Ru4MlDKmWWtxL1QmmU+RC4avxDUEUHK8oUDqJi50LhKbCM
vru+od1vlsu/0qvo4LUZs69hU6fuSan+6jXqq1FChPMEugVGpYlBuadOX8RGWfxRXypHIwb7IPcP
Jq0RBeYTEd/ReVoj/kOR9K25cSdCnK2aK+G3xXRxBFf+ZWKTbhtMMddokkZs2ahpRp7pcDVDVzyI
M2zG6Ew2TC53fF2Hjx5bDQYrjDwSZIx4ZV1zN8+Xp05duPMSXIB1GLe7FPDL7J33bgku2Ac4Y/yq
d0F7xMeviu2DRT7rUE4z0+X/IBBDzh4+t5pPNzcCA0JQCepSPlRHNqm18gOPxsfLrGB6EfbiX+ni
CxwN0NHlht3hSSWfdo26Mcveoq+ChwQtnxz2ha2keEXyQg2sgHuUF5hC3Sw4OEqPC3nTZY0KG9sX
QRoGT6eJBSoWg98lJOWz16bMeG+Yo8o6MAUlXS0fCTmXLxMu5FHMZCVBsD9o6ttXjkLNjFZRsI9D
IK/nu/bnTxX4a9aqrbjJSeQd/iKsEmvKiD7AW3/AmDc1WEyhZA2N/9JYeloE0YHEnc0mFqMpwVpg
k+1xyiVZUjtiEf+uA0WAtYRfDXq4XSdUwoVmtQCvi49rXONDZulYLnqnqONPIv3B04hGdq5b/FaI
Ju0LZB9GPkwePxEQvC2B83ORtwRWxTMGpnehKhDbwwItiMVdOoQ/FgJZTLfGO5LgdSspyDa7g4wI
anqwwwOE+Jpsm1uvGTNs/gEG9y6+SNzE6dWSoM6M1B+RwfMPeecdU+wvEpoJmQIF/G1k0fxAs7+n
K4mDn0GmCdHqZZ6eUFX1FVKJkuhsghx0FcpYBFl9SZJcRknkOUNeX6H3AdHzJSa1SIPBb/qNgZnq
upQ9rFMHXWe4s4rB4kk1j4RzK+diOvK/tEsHDpqXrNQE2zsAkjGzOMgE510UFurxuoCMLmxN7qFA
TZidyZ9jovMbiDZJNpc+bzKcRAxgom2/Q7gT5ypXqCVr/DGAlpNxoxtPacLRWRruuS3H2Ri7CGnT
frIfDbh6poCkSbzRwib310Kftn44KQpr8oKBWmhyRdE8fTKArXg6sDv3cHjgmGktrvXcQvhgOeB1
/BI0CBdcRkDMaujtpYTDiUNQF1txuxae72QBZJ0qpbehqzspZIPwRG9xMigOOQ5JlLOlIZB/7DHw
eEq0ivGuJelCxIXZLQQCSkYYRLV/rNuv/bbdaF1Q3X0xh2QRsWS6fIS4/KHkba/lExh3cKzRXEbl
Euf/N16ZeePbwEZi3fdi5LXTW/oXblKjH1r2zllYhFYoFtQy2yiz7gytmU7vLpKJJoC8Ae4MGjj3
qJUppsRSd6g62opkan/8xiivDef6hXRxr9DzAMoFvlZnB5ZsUsNNvKAUM36AdoWhv1qIt6wKuhwn
6AMxLj6QBCnPXQYlAKRDQoUDb0+7DaRv6o4J4MzjEnAS0ELkpU6iwtUD30Ym6Zyqi9LkvOw8IssZ
JHTCBP46wW/DduPjChhKLGv1GHZgsipz9UwmEmqLS7xZJHnxwLpYhGki1lbG3M9ZoW+54AZd9cxE
mMiDXy0NN77r+uSot0frA3W5eEkifh5+WbC99fFsuMCaR0KOR5zgGzolLYDPWz+4rUw+rLyS9SkM
n858RkPDkCjJUfBHVP/fUBs7Up8k+JB/FRIM8pQxDceOFnMouR1IK1N+evtt1SXLRZsS0CwREtzZ
Oh35bFNMFxQKJKutvD0+d2wobwtLx4x2SXlCGRlCmlQzxWOReM/jwxo4SnLGxbJ+9JLGm37VsuA2
NC1N3Z42RNk/l64HWz6KSvk+h4MsKrjQiBDfEupLo3yTCeXTNW3eA1I8exPh5981WrN5n5J3iL6K
JjGzHjbA6iVCxuiak0oAuzkyhTjowj/9nXfZhtFt5dE+zFG1N2i6bVt2SEUciqAIsdnn+i2A7zF0
2kXOhCEA4wRnVaNEsCkrK+hUYPwm6QDs/79wPydKsItk2joVpJJTknQnKIGoJw04p0pQ5n1FqIb8
92MCTqQdSlZP3J+40HjitcOJDpaA4Vbo/RW43M3rZeLsHx6NJBuVujPQiDKzxATLJtXod2udAbYD
wETohuQtofICK0LrthishPFJ7yfvQjynutlIuWjcq31OiwXt62ifwanHauXq/Eqp23e1YoF4gm6n
jhHnBCnWbpp/qR3b8oQBJjZfnPtDFlhF2JPeZDrgNdPyA0X8SPkcxUas6F/w/lCpSkVUyaCJAgz8
c75zi6tjabV891DAETbDCLz0/3jarrJYYZD/Wdtkmugf3gt/sva5qTgZefGO3H6nDOzdqQHlVlm3
w+LHm7/2VWnsupgQoZURNA+6AMkf/3b6qaEa1QICYDjCZOxJ+Rz4ME26eyiC31W2YgxBZrmVrA6B
r+NRocZhHumqZEPtWYjs/C/cpGB2/7T2VlDaPK05wxO6jSlfRd/LpnAEQAXULT0zOGbDyDRuaf9z
4nl+AObCHKJ8ZOOAPRc6ZlwvpRd/rBMawFXD7oLZ93haL1xqCWXDe82JP11R9gGUXRKTI0CHFJ8+
G2X+ySDJGI8VCvYZ7nEpAO3axq1rGbEGIrsx1ZNhzjzF3hvWTXsX9a09I4SvU6TkQn/H5eFmWMvW
kjFfDdVi5pmex41Aev1MI6Jn5R/im8+Gvg0or0dq5EEnfYXu9u0946MKiTcfneSHvolk2j9TMmyo
32sMQ9iuHKBnH1LuMPp/zpr6HezyDPICqRqN9sNA8T88M/y86dK5KbO0PGehcuo0hpXw6rCqBvNP
UsAT8x2HmNZge1tDzLoX2T7CN4BH/gZa6Atxcis4hnkeNEIghwjIUI2tFf635xuF/8u9D/kT/kt3
vIlRiR+M1HqyyxdLt+jGT4Ip8DopxB2iwneIsYztsiFbnt/EXqVnhrSFuVRJMSBUKsQCGcObhMm4
adH40h3LZbe+7/pMx9ANODOHeacbTTd5MGy2TtBmVJ4LJtUOEVHq4BXF042di2q0lsQu8cEarZAE
dIXO00sISyb0xKKipCAYx4R+sdVFamEbK8A+15nA6MW4R6Hz/jzWXdbvWXGd3nTQoj2+BQIssLXT
OXpXmELPt8jMouPCkdVIJJombP9u1RhqUtP0fqO5NCZNtEC3E9gu83akMdMJmpLAz0+c/gOGur6Z
A6RSrMXI2OYmqjuw0g7IQ75gT1bhWKTfuV8+/7kNaF3eW7R9hAMtX7kccSvUPsVPmElPRQgHPVeo
nyvXwaw34iljNYTkVXefHAVG7zKikkD+0IyccrjLGeKhNFNvDKVFP+YzMzWHHMP+QVHs7b5HhxFd
7D0WENdZMiXacV0h/ybpmEtHwee7aC4DA/LJK386hcBVCXT3uQzj81WToCVXtuAlxDYkF5iL4C2w
KLplpDxUhiTZ8/2cqqumoZbUQd+raAgbEnGbipVZMLpMKNL0x2gX0wvcTxf8+jrFux7gDD9k7EXM
xqANRfZQO3+hY8C6oSCVaE1fEje6EUZ2qCdZeBscXsGUWhQfrBY5gKczqPt4X8jnUYQMhHZKL8Xh
egnQgx6fSIEFaRxxsKidaBxm9Z4W+RmtydfXWFRpD2C9mINo5LiUBhJ6r1HhVw1wYvIMMPWLfPX/
loaoikliqhPgMVkiacuvkkab6G+7cpcNh+uH88sIbrjbA2oYEQ0FMhIHE7IRjgUmE9qmeepa7iS+
tkW0pT1e4WnycL/fzu16coMbS0cBGXoAv1GayglAS1Tk2siuy2wrSNzin83AO2+1+iPsprBSczIo
vd+eHQWosvPw0DozCtDefgnIGkHY2Hs+0h3FaEzwZNhSew4m3tlY+UYcT0aN/RNiP7MckHKCBgsO
y/Y//xRm1ggkmMZ5OMX9JO2H4lZyioh7I944rGf/L8pvuR2XslBxFaix94ly/LeSETCbq5lbWd6r
Q9WN8YrcoPZUsty3vylX8dYOSzQytXEkgQ7xsz7WQRKQjwkYR2iv4r1/1DHAWx79zCC+mZcOr0xk
9lPeTrrs4j7gbjfWmyuhcgouaWKs9HezJOqHBXfrUkTv55OwggI7iy1aTxvdX91VEbUozvdxPipL
CjSXigpUyBimRPLu5irEUskSSqAlY1wQ8RRt2ERa+E3NhuNs0g5RWY06Ds4x5aHP7bCTYt5Q4S/E
DS2EMdCpVeFeB8NSdlnLqEPf6YrN3y0Eh7MXuUYj61CUHweFeMkYl9jpZUJWSg2LCuJNmsf0ywYD
m8tafkhDOAXf/3uBywmJgOv3ubmlQ+r4tzaQwOs2GxXkSNT9sw0ZToXTLZpDoMetAItMU1Xj+34u
bA+ZpMYdaX+iLQfXVwRBLHvamSETCY+FBjxOnZ/BH/v2vS4foZFknidyZGdm+yI5zRoNAEKlrYcV
bkBa3vxdZaB+6Y0MppLfHADITTvKO3JghOSmVlpfd47lZZRhOxd/YJqeWmfZM3bdxS9FhXm15RML
cUvFD5xe10dVRIPYfGZb1oqOSqIcjU7EnomBFEbHjKFJq9RGyeoSR69AyqOPpcOTUt4L5ECxNE6T
VNDh5TMA5hL+7CK+3pmeXOloK4i439Tn3qW3UMldZ9TE4LQhWwxgANZZIDsEPoLVRV+pkIxGyRQQ
tQzg8YNTH4aLHpqdaiprPkhO5H/Q11uvZv60T1hXVOC7GMB9s9670WLgE2Fai3dwOJ6g5SA6liJc
5uomrHqq2IPFMlliZx/0MFbTUfJNkcW5wjmnODdvUVVkyV+qzujXuhwdTrPdg03mEDWbCkPlFqkw
DVwPnrM1wgyJO0BMJZLHomoP/39WPbER92Xfu+hY8rtrbntXHNRV1ZA5+0uMn9BKNynYdS+DK3GV
IeFUUb6MOUta1UKrJUh13MjNMe0cqr/YnD0tf3L87fsOLpA1If5o/Oy5w4a+yZ2J1FtsaJ4Egm6H
1YztGgyOdY5pfpqSBCHpXti/+r8AAxRg0cnuZJpQe4kWeVDn5zQdlm0jn1vqCpnCTFXNeUo/zgSM
NGeXqmb2uKTIv5yA38pS8mRWHg9qEJ9EnvWUUD3DqjCPkvmdxL0hZm1D5WATejYR4wG5n+B55oib
Qq+TNxGpm8P4a9kMF+RA5l3YFa43Y9FFxb58ltY0AhB3osUHD2wXerjhLJ4IhKJrfLcJtB6G/OXw
ykRFQZqvP6TQ44Gc73vrjWW3Ewk45MzVWUPwOk2IdOP0b819Bba1tOeGpUyLaAJNZHiMEsxNFgF8
AkGY+WPphoZH52H7vAmxUmfCAxDDPv20EDXxTKnEnmeKAg7K/2WUjPBuUcPaVSCDAFPGT44ajjdn
X4jynEbhcODaAojA4BNJvQSQF5uQV+O6TqFi/TpUXd87tsO+Pw5Yvd0CslkhpCNrWkThIoZA0h37
Gtfl0i7Qj7FSrUiNZ43zIdqbeHlzfen2yLon76aKbl9snquHJyrFw/yt+NquKc/egCBd4p+RffG/
Z6NVLdShszNjJdGkTbHvCganrVQpJ7mDbBCTddrA66wCAqw6WnYqXik1hFPPqldzzI+5NJmne/E6
yIg+5lEi6Q3/T7PynHQzbHUt9TbfA9E7WLn4dZGnTQ79skWSm6HXSUlOFziCPlPARdUaM53Hb/oX
ZvvWjE7q79Sfo4akPiJFD7TZKK1RxpMNT8X4tiIq8nENRVchPl1h6umtL/MsbLayqFHyvQesSRVy
obRKxOUG+qOedjS97C2sX8+nrcCIZETKrYqkVZZ56cW5DMeRNPFPfsX30zF7OvPFf2Hnv5lyLNsE
qVyD6hUacgv5aSmR8TrsESPz5B+Xk3CWNN0z6Z+9za21uxwTA92c0XEgRUlOBxZ9W1ehdxpuewyI
B+5wI7pQ83J2VVcJ+Uk/B5LqDOJ4L7H/USQfW9Cj/W8bP4GMmIs3vm7O/a9mChvvUlA9RALYNChT
h8ndoo2hZkzTmQwTx2Ws9g+Q9VYbFT+dJiYiEIFN72PuHnjQU7J909dwLCH6x46niwqPO0p4Th9+
5MpvtnQakAWniuhNSaXkGlC0b50M5wmSUMzPUqvdm8H6Nwsad+Hodx2SRsmbvRV95hA1daGTPa9O
GQyN6H++sPEApIbMvWCHFmtxTRdStxzyT6A/UDImoU/UK6RlWlpVfw95KkQr03oQzr3uOw5PW+fd
9qt7nnapPoALZH16ZUf2re+ZgMmnBmJTZP1GU0fSeX8GyyvOn3JxOzChOvAXNsezeghKJ6LT03m1
QlRTHobJPhYoMK1hq3Bfq3l60p/09Lm3ZLsBgRMSR2XqDef5mFOf2kU5xb0WvaS6yvokaMFGvOXE
vJ4oasGS00gTJzK+G5qoiJfdGyrO8HYd+8j7STarUeyLcULHD1tmqVRT8xf+hNet3NJcrkmsss0m
O0IzYRlrO7XOg+x5RdSo2eLBv3o67kC/t2Qz32EwXwMSlLK87yzhqq8aExepqi14GdO5GEapjlf9
Kw9iY7nLhHWZbafWXaWdfk4/cNSbxYmfoWAkbF554hXmolPkdZP+5rkvw8YJCkHDltI8yN1MoDms
vNFF40nK/LmFNRgVtCBVDIsICKmKjdq4+MTntF7XETCaleCj3I15DNppSofd0/sHaEUwgZ0zET8u
f5v9BFGtCJCKa3i3y5Wix4XrWCSN2DogDZYcMUPNzjmVI0nRMVt5z2vfmz6kcP5N+1C17II40EDc
kRCjX6vPEpvtAtPH2f22/0KZeFjy068+rP8cj1zi3r7AEZWDgbTlIksb1Jpj+xgWUID0E4HWs6+o
+s65ou/rwOLkYmVmFZkUEPMZMVOMhYQi2cvjULza/FEe2jjHJLQj30+Wt1MwDpDwIppdvEi6ORca
56ROwjRrQhbip83OdC50hf2YrTokMBV+7TI74ZKTJ7+Z7o1ZPA5/R/oNO50cwz2Vs7MvxITPULNS
6kfcPxmndx8lTSWgbRAEt05zIdF8ryJrWmoZZjotOHoMV2gabiOWAhvIiJF15rX6vPhTl/eVzfEF
3EEZbW9u652iDtqQ9Fzz316si+gaGo8Hx7kFNvq0GMHbLaNJ/HxJJrzMtBQ6zYFeqtNaxz6XgSrx
raQFp+YzYt390ei3UdGM87JuB4bx3Xc7Fj0szA/czf6XCn5E5WF1mNIT7a/HL2xvJz2ghJEHBmd9
x1lc6pNt3wuV+6anFW878pq2uhyrB/lTEnpMz1uVEz5+9hdJhMaYvaqi0Hy+OYzjzFvQCdJJNTbz
ScOOHqIr+g3DnW0pu3z5LiDi8DcfwS7ld2zxK4bQtFgOODkbeDxXGwJxhxq9kcI9VWmKwkjmPVtC
hL4vb5aCAPk/DnpC2eIqOIhpzSUGQJzXHNEj2FN/VHA7Gjw0ro4gkFkCweQfuDJOshDNLuuSwR0j
AaXuDiGdM7u8/gV0oeswhzIsSToL/37ouTjTEH5/j/kq9UzLtAcoLc5qvXU9oa+hKhBOgAJ1pgpv
ToaMfzoFLb0NYP1ILckXwTRWVpNuppfovjOB5R1SKNyfLVZn08qAB9oCour9EVxkRc/cJTUtnUkE
4RjhX2ALoSSozCPaGwL9zGGvlUaFVTLol4AlUGsXHP9BntlA3f3SLKo1WUYnnb+6UYoODHXgI7Cx
pEpDDgGhzjg4Pcp+/Dx4Mnw03Pz3skoqIzB0YSu5/cbxaevZnholR/IaevKFItmxSU1MaUJ4qAb4
gQ4AZv+YUERTc0EPsnQq34mo5MtLmEjZ6gZZ/BbJPwefGshW4DPzwl5Z1ZirfJYVgevGl3aU2qah
u/so6Et6LaYZvlpL1ALpTuxVmh6L98aV3HjToLmSqqjFBkj9JfL1fFVAwcwuwOkNjVo9BY/Cwup6
ZMbuYdQ9XT44W8sa1xq296F8fJmODavaQEmEwnmx57l2sGrPhXSC8m5pZ41MsR2NOnHvzvzZq3DI
1/yIz5gKw72FZV6PY3Bn6scnBUqrBnn7FgSMZwwlx++AudvB46sQid1CK3CRMRYLbpnxJyJXqXCp
DvxiMJ6uXvTHMTmmS3HIR+fMBaircfRD3d5fEKQPO4e2Jgy07rooeQBjxQ+qkhocJfFclkBNkTXe
hZO7z7jwx0j0rIC1TKtGKXxaeYt4BNQyd9VvrvTkjHUtGLvnR2ax5BMxwWyDqCZgI0iYlvWchRqF
tej3pC9ucGMTDj0TRIeJ0I/PbD01EaOzQnD5YB8CiABsICTNNrlAuU2hHCX96DnmtQGznaQAGadH
NJAoyMxg6CKZq/TUmD26ci3OYc2h4AQO2jiWCJKKBHqzhCG78nbQv/ac5GceU9mbhzZgSEbwgTJP
rvV7maB1MFwt/NYlpRzioJESZa1b1J03udi5hHRVmGzojjtMvbyrIRiQ0M+EML109ZvMPd2HDBRn
A11wzQxrl1beL9gNJ8MY5bfRYbDq72o2cBa/2C1B87DQT5K7RqmuKZhslYUrIw5cF+L16T/ZS+95
0qAMbfAnmS2Ir/i5yxZrgANLSsO0DkI86O/9Zfh27apBE+9CFqOMW4tR4Zq2GOPfgm+dcDYHXy9F
Mz/LN7YPzlOZENjpxOFkKq1Nw6shQYwSjgAHGNWGCkX3PQDBjlLFxb0gaW7sp4mwXLn1GGAv7dl3
VTNlUksNR9Z0jAEm34+XTJRSIVsVsuExnTNjbzu0JCnrlqpO4qNPznmP5KkPbSIT3FTy2L+S2D7v
kiNDYcbWWKrPbzkihMsYXcaPu5paZP7VEaKcZWHrkMjpeuzfeDmO1SqgV6vaeB/+YmNNYEQRtpZx
uFJKz2NgF8ybZ2a8bSbPCqfXjRODkAJGipYU/HyuCwHqQ0qPD/2ae/zQcnESe1hvsH6AHcLnID2P
XM9P1SexSL6Rt0q80GsJJLCkaNwlA8tJt4/iVypeT3nIbTJOvgAaV4x06Cdhi4sBnpAsgSajj0pA
9jsVgY4Nt0HPIx4yHsNPdBJr2eCcZLzgVwhYx6tmoXAVm51WnbaO3grGEDhl7aO39bWM0WhQkHhQ
Sgdsqw8T+Q5T+HWwhZdNlLpjxePJNcMiRX65jT1zZJ7x9oK6mQqBauk2OSaX/ahi+TZTCQRZ7MTa
6s75k85umKtGTmCDIBcePAIS8PB2pgpf+K+1zmmM0DAxs79AkjMsHRipX8u9uZEhIQqulpDzsCsA
ETd/+HPfV43Id/82VnITdQ/mmI30JVU0gzy6cBcseKdBpVtQV0gX04OPR5dfnNdpOJBjHSjaVoy6
fGdsqQguCLMpz9gi03Whg3KDu6MlouSPrUFqg/7qY8yMXdUd4qNo0zjb9YtQ58vhCTuzr+HFi1il
KGvox0boqjCmthhiDYaerQD77QpioKfSrE9yIk/ylmolKU9nDcqmVNi8OS10Lim8uSxf/i81ci2S
GH2XqrdWGX78287n13hiyUK238P0DPhONATkFK6GKwurAxGZ/9XkJDQk6O2omLwmzQ3YIGnGmklH
gDqgpanGNOBvfYeNyUXIHgey1vfUaNsJWerDfe+RX/p8ZzbuSGzX+h4q1i5NBqq5rFNiX5U8hvII
Fjha6B31gF0AFcJGK8awMjJcsDpLtHpdaj1RppqNzeQjvEARMk7Rv5Wv4QSJo/AOT7mIr4HfVzBT
5HRF8Uj/Z8OKKoOtZHdDFXbeqmUwgj9IHSz1abNeCsa81m7gL6r/unQ4MPZLzUvLNwK+RT+XMZPt
4w0tndI/UQhjJXsjXv6+GNgwIfiVZGVior0FRihhlMN3aXHaOR/lJt9cG0fv0j+sBUNy+VbbzMJO
SydRlg4tDjIMM4+fU44wXNpuMYN5UznEJVs7ZCWhcHZ8F4CVJhOBDtmoGygAReju+KOWtWEmPAWm
7nM1czHqwWHBtzGtt1fDqHbY2S5FKHb2B9QuGgkQCIFrusMWVycmPPk+zPJ2UhWBVHvt2KScO3PJ
flzaArJspG9+8FkR/sOJ56+LGccUAkGS9/vE3O+EWYAyPFqF8N4jf+dzfIZyQ8gdth1Bnv9WSw2S
puBuwW6QcO6qL+04vQQ6aUgUD3llabP6ADb2lVvAmYKrZ8787adVjmKjlaXxEtFLyQ76jX5iVrfP
gI0L1cUQg3Mi53bJgM/jPi/omGHpcuSQwogRo1OddOggFqCZQEBblEPi+opMBOv79xIlQ9Q6+S15
LlstcibpLqa5NbC4ezG8fE6eaoQhQHFS7z2AMCR9WFgDbiNY5fIqSIf/rbOYqxNZOo04d8BZjZc7
Cyza5G4XUTXzLIjMNanaQ++e7MuhFyFJph3126Og++E4UkeqBGGiXfkNNLY0s7HZW3TsGI9lkjWF
TaQL1KBRDGD6wBGGaN+rUivo0H75hfrXDidmZFQMvUUxa2+xWcStPLr+pzUdFwD16RxIFsIn9L7b
s8kA35kKyZdAHdhW8niYzaG5k00/U6Bh9mqxV+ZssQ0maV93FQhb2kSSoVQHggSg1ogfm0MBPa+A
fSvf/8nj/JK58IjivvNbji7TsaWTHa7Cyir69umf3Fol1y061WyaDdGwZEz4Apv0ZVPPYRH/kx5+
A+o9iifkZBYoPh5qofj1aXRttcSPMYS55TaiqNa4d8gK+rmfQHcivc1Fr79/ufjlwxQS3o0CriP/
E77zrLvuuWwlnMbZ5ZGjzbdKEBYtuYKbt/RMXm7Lrw7367RTUSVkoDeEN6FOTM4+EdozeOvnejcq
2bVGE5NrNfa+d4wtfNZE/v8SP2twPzKZKzU69eGwH7nIINu/DTnwXX6dG0zxZ9b/1BIfi6KNqbmw
EKpqc9MDdF16BnYMh0a0+2iSaLbz9+z9JGWz12Z9n8dfaZv2y08vHkncK381Rlg1Z+cWlkUw1JyV
ZkdUg7505awa3iwtTSFlNL6L7VjhYkfs2xbGij8XpBeBeor/Vhp77qSJi/BZHNL0DbTys7gr97Gp
t/GVqVRUWTtu17pREfybOsR7b93tulp61hGnuxBEE7bld7gK6OGeEElzM7rqlhinJW040pIfd+DV
LizmcAeFqYduTFFP5bLV8+kBAqqD0yR7g16m1W2eF7Azy5s0LtpMvBgKFatDSUQw8dbNHWzR+SGM
RYTSzZxXQeqYVGfaRgqFBVuQdz1hhwNboMzj3QGcc1+54BZlk2OR4LNTgXrjF2nyAuE9PPM8ogkG
Ktstb5h7ZQtSOFocCIeMBaQc4AqHZ0lhhBPtI4vnkUh7LqYEkesZX7KHLhFeDREBVhsIH7SqCdg/
Gaqny0Niro3h2SPZUgf2ky0KAFF1wdc9PGfVd9lF3R3hTRTohNnhGOKTxRH8HBjxCB5aOCUljEiL
tUGBwa3+THOhE48WmxbYMT+5Z6aCp9TrS5kf5BFjHuQ0ft9QB1zYXrcynGNCPUr5DoYMuULujthZ
USruWISR+dm/tuSM3nRkKt251A7j1LshLkxq+hVuMxZpdRjixeLfoKTvB/uqp2b6r8dgSR+2GO0S
tdOp3VVhGejLvWq3rnbLV0P48AQ49Vw6jjMCQlA6Zj6WVbYaFEEfGVrPBKo7W+N3mEFY8DP1ry93
lWNk7OEYwFD2pKBvIfYizKpMSfEKDKG/0jPheTLRE3eGdBLcgowEQ1vEPaqbX0B7qCQdCxRT01Ru
FEJ2fOft9qJREK/YSN7SwiBzbDkQg9859xBTzcopdivbdJ5rrh/odODV6B7oeyYVu+ZPcJJm+AVK
bzpNxfRbL8eO3Oqk1eLhjcq9JG23XyiOMvsgWOejEJL/LkQ9fxhJFOxzrYLi2It0RFn3tpjhgC+G
L/fHx7WIdFH06LlHia24iX62BhxJXpmxTeJxhOe4Fo/W0mYcPby8FjNnfBxi0wUN6m53cdYzXlS5
G/5YIpSFtqgxGHCLW0vcp4iTbRToqWGpZOPyBRrIWRd1t/bdgTKfowopCRX89TZeIYDJe3hLmvH6
4E8Kh9zX+2nE6xu1YAJtlvprc/lkIB/blMPnRJvecWTypkyYBP+QyYx5SeFhVt/C+s1O5dWjHg5v
oxqFIc1tSPsXXUDWSjHk0+uZs7HorxjuQn8nymyHLiz6jndUIdUIxRhirm/Rl5RAOnve3qZbx7kK
gJzu5PrREI2kwXLj8ZdOGNH91x7iDMywREi9GHdjXIg2q4N21Kn1IRiU7S0zas+mOgbd7pZitx5N
CBkNBbbQO1WPY0fsCMR8Aa8UdbwzSgS9d65dWfTXJaZEMH0PBtjTi0SHuG0mt010kMBWKwrje/eR
kH75tWsmUvTF0Hn/pZq1B9xi6aaDmXLUCzS1nNpk/W7mqcz35vOXshnCOyFIcsIy8lWmwPJig6eH
iXiNvvHFGrRXlHkmoaUNy04rUcOKAAG0odI0PjNvQZll5Hbh8qISRD4dQLo8J0zPMyhIVPE9romb
YV2P56jMWOqhMzgt+70Iikfz7gXWw9hqXlRE2LBM3S/L+11ubwoWekSeWRUs7rimMBWHgZzIuKvt
DapRQca0q/XI3no90vH+TElSJ7m96AFJVG8WwFOK/HSdsufu75gpqALkleJNQxhQY6XlAn9rfus3
khRqdS/3ujsfkkfTBxvXswJCkB8h3yc8Da9x8f4xZjPT/grKvXZUf1cDrqcwYO2NdjQTCmIyDhIO
bVZOcmaGzALWJ1W39s/EHzQ6JBP3em0vHl+HAk29m5eKlpGb1M12TwxSUnSg9+7DKTvqoOaqqsxS
vacMdEh7xP3k1tXvUJtImYyrdDlK8dNnMDDgNCSL/346+AMqwBZ4K+Q2eTdyHP7myODcPwNVfxLQ
rgUDuaMiQ+ypoHM14YDqX2kJgSJaQQgnSuqMGW5ADm4t3R1RKe24CbRKy5CCSAQWnwFPOh1ecpr3
Uv4foayZ/GUpjH24ARzbDpZC3A44Oym7Zm2luNJS5rUJ79wZ9knK03rJ1xnHEvljDoJxyGlrobYK
hw6dF+aXIQ7IFNJpMeo0EztMBWylIkrrn6X1+mkINv1Ygn7SFIcSqTlfvT9FH+Hr+btFyw//jXfY
qOgeQE9pnijZuCM+pjehGlXJALE8ZtoBlHzrZ6lL5PfAVVjltjvLFFwPaZrJQTtZ3oHp2uPDd/ZK
2vl9M0kERYEzoKnG9vtWhZa6yzDPoVxUU4AFD7JPHIRmCLvou4MtqzK/uFy62sX4rt6sNMmRq/cu
s3t7E64mrp5QKkddAlvfrsQSSXd6N2B1woLN4uS9q6GIMmOXjF4fhdGOyf2A0sxpK3z2TyEBwMJR
8JAdH+sq+p/DKeI8b6LNFDkJdU1nzRtYU4jsy3lkoKF3hfHZOLnaAYtKc1FvCrf6yceJ7NEC12BO
KCB0uTr1cJaDCx2D7TeWo6cHglwJ8dszG5+VChtJfeXkq8jjsRY6K9jI6e7iiXSmHCXpENyUIur5
YNRwMatBvGDQYpz0p33vv4M5+8vDGAdoW+00sRsp9CsmBgvlx6f1cBTuR6azV2GK6xGLFRA81JfV
HcpHlEc2ziTBkmRDhrRGtaEjPhdGN2YOr8ADPdXfAEk6N9Q+XuVXloy57VBwbOVI3ciO1Y8fpLXP
vfANet+YxoSsT9so0J9Zc0u8wWHyWCo8xnpxAu35ImNstD3pM/aUlxVKwG2pQDTSHIdtvmcimHzp
310hc3wpbP3Drdpu7HAKQ5A2rpd9xXwuI7vzzWExNUMgW5dIQHRhh/Ra3zPswbPmVhoIr4rTY5hp
0PrZejQJwUM4PufF0KyscK9B6PhFZe+Yz2DCmZyl1M3ZLMqr25Py0zBaVP8HQd2XAn2pRKH1NjQ8
qJVNewxRY2G5pnqqgDc0MWlBUc1f9QwhI1Ud5FfD+CfX9ID/dndUygmwmAOyXeDoKm/mO8ikF34O
P1ZVbnQonFXA4BGo88zSJ070T4lapqo2QFa8NsnbzSDlGqOm1Y1L9V/GJGasUWklo2xj+189A/FY
0zykUOySKSnhM8iJiEU99LKUidw0tv7zz0BXocxxDtPQShoqEd7N0ZHEajnHTnnEsalaHRNlzzy6
LNNFjvWFvMqYaJLiw4CPSizXOVlulIPl83lSmFwXSWQWR1Yot5bZ5egW9AURk5dj3DfQWd/1DB5s
IfhCDke2aKat8o7HvXZfAJVay3ppN3Ea7xp6CvpBDyOXhSDfb3xKZcPxLqn0Oa2LjB1UamE8dGtZ
Qm8Q66jFICl1y19myo1LASCU1TWvyk0PJzrfnqtP5sdL9sh/MFR5yD3Hh/C07XaVaIra5kIcoMF1
SsFzCeo8yItpuk1LQER7JCID2c0srfnQ7HdkJ33ulKDFypstmiz4AAv+0Jz4MK9GCA3lLmIEqueD
TmKEariLxkUuC8kEjzJR6uKDgk9ZMOmt6GPQ2nziki7q2PwnGtcFeNoM8Ep11U/ODwsEOX5aCd12
55dl4yRjZ1bHfaiipZmuI2z6DGu5JeXW8BXnChvXCHVASzjjpELL/rZ7Bi45kVgFtEEhmLx4LEQM
e85m5Ge1XTjyk3oXNbv6/7ifF22O1hNvTB+QzLJuYaXxckUKtzGQfsc0jHtUxX0/Hq05MOpG99iG
bg3t7FepUGuVN+oLIlmHe28PsmGzL59GqtdaiZaamWR1iIcom83pc20n6bu7IZKuXDkgb1V9xuUI
cXKUK7ikGqHiHKXN2EryLA4oFkrpUFm3/i/9M+KKk0x7IQf7XpHj+g3hRps7pcHIrLUkKMgpWz0g
qBdsUIoylVBs1snsd18tHex4dbhg38/WLQdrMJXcZEj0oyGlP+B7D+uPP3NFmWNazSrQtewKVZ1i
JG0KQQLndctuC0NJ18LhmNbs3OB1lNC/Czqn05tDVHyiNm980W+9uCAX2V70tvqTc3eVpz0ZU0wL
dEYW+E7Np+F1PJQY2ksNUyXtAdBEewQXwLVaIYCkqpDkyuSAYs3FZ1uGXID/bY1SCJR9MLY8mwfJ
CwkqProcvLHZbaq9ljiJ/gcCWacUK4HzMk/QdJwy5PelE186uGlaZDU6tKAxixF0evIvj11l4PsR
HjOCmX7Q9p8heQvMT8FQrHlSd93SG5AhN4mpdgQAzWSKe87/oZZNsnoqzd2Br0BeuS4wQpKLZagk
yJFLjx08/We0wSCBl5ifGj8tIFirhqGNp+7FTOZFnUQMgziwA8nQjnyEoZbFoLYUUzkaRKOL9oEf
NfdQUtNDaNnlVkeLRMYB7N+sK85ATAuCSPul3xalQjSy7RetsL0oRHvITjsa3XAPQ0E0eH86S7Az
qbVsL00Ccwd/lLpqQYcrhQSiY/1KZ9PZPB/cFr0r6Jq61gAFNB5gXeWpmMmXfqyRIJBSILG1ekbW
1Py0hCFsb0HofBr4c8VveSLMD+TB7t56N+PA6U7n3jvrleMTGJHoYaUvOJTlrpy3T5rdBsIGenEg
A78Kl2BonzAzTQ3LrGgX9Ajn4eYSh1teR7U74Ya2MCK0ybqEm2Rsxqr3mJ4qArUhSpjZ4IkmN7xb
h0aP5yeg0WMt688QxmGUPHvhjZBH7/H7WKBW9Hfkgr+RkWKwRyj7dCEePwueAqzr+yZ2l8WZl//x
SS3m9s/N3AGmPEOKWSlFzlG6UErG6p5I8c5lE384z+OiUqZ/sqGKt8PVjr9msQ06/ZDaGhf2LN+U
VGPv37v3fBP/2O4a/jLY8odMFYlke1p6seHL+xIWaiWa9MXMKQ1ZB5tpr/h+tgn8UR+spewHh8TB
OkAunUFkVIhWqRBMR2A5+6TsN0u006RzkfCM3TDVChoD62MwmvnWR7bQNqITrHrSllDb18Nh9fQ/
1ZFYoU/tmut8oY8SHDh22vxn5xQdzhFixb5n8wmeRpqTG43H46m4DDrOH2HEFufGe09XdJdZtXdI
hDDL8CCjyoB2elTMjYBABW35J1FUnygr5W9d3iBNa+LH0cStTsNSfIWLOo5+TpvU3U0S8+hHFOtu
HEY2E/MKKSxD2PhGBIaWHvY/MFJ4vTg2EyVuhIQUMvoLc/32omkNZWhl5QBCihNf0yrBfyZoe+Cv
GRkGyv40rpzN0nL4BJiN7nmvWIQTZ8NlB++FJGIEboNvSsWGDhaelO/1y5XpXvT3fTz6hfUEBu2z
VSbf3GTxfy/n7O36WT1XY93ulQNKSKtJ4qLVPeBIycBlXD5qdYT16Dlci4+LTekdH5uSjmgqyYWo
3pZ6JWohhgMcarYaJFgGoI68D8U0WK7soiVXmomZunlzQcPDRmJgqWSFKfo4FnomKFZinMR8Ry1Z
WDR+9HhQw8+3qOdznD3SXqZbKUAYFAVsAyhqJsaX9osklJJ4xcprIMvRMPRI/ZWwScPcdvJC3gSx
TAl4EVD/VRPc6RuOkKL89CBYnsaQCBkcBt9ySQjFzBlfXl3VQ37EjLn11k4LJWlbeSUXJHobw/j/
cTvn43BeE3kLbgkE8WETW7/z+M+UJhGq7maxBZeKo041+T8syJoEuAZ5qsK9Zk4IUxuPwB3HfdrQ
hI0Lmxz/BOqsfUy6Wk3jkgt/JhgrYGIklw8XT8UvADoybv43pDrX7YBuLfGJ5srtmNEKcXR3YShK
v2yl7hQNRlJuJm9JNXvFaQX+r/8YyiSBG/fSt0IuEuYm+2jC3vF2IK5vQG7ujfDz1vav++aFuj1c
z0Nx0w3mQmx/vHTqtauc8gtjehQSWGbxMM5mAyvEhDZ9T1D5HwhHYM0kYovYqpu4mZ1pzaMu4+dF
af2Orp2fEE6Nr1LbnYSPjd7pBZeP/uiAOZ+5L9v2iR/wiQpR6GiTy/DuGbhCWnFrfI4ktJFxU5uf
0tNWG5HGAkc2jIQcmJkk0+Z8O56Y2GI7EYFAV2lE73Zy2d6jklThAL2XV9RRHQ9Hmr8iH+wLLD8Y
x02ZkER1i4OMn90YTrOOKeikQ3sNwyjfqInEowKXm0z1LCoKyMeHZlrtbUuGf0rpx05do6ohTGVM
OEZmc79fj0SWXUba4bhPqBY4XN0I2GnLyVQee9kZZ54n9AB5WUjeiXg09Q0VHFjh3b2Q1ZpZvZ+d
P5FWbeitWD/n5qhiSrlsBhFeRgAoRnoEXy4c++S4vDOOko4ciC1kJ8ooyeva+15N5+H0I5b8NmZK
EQzqlQX3z5fdA42LiyZhHNVIu9+MbcnmlR1lIIiPzouGklimnt3RQcd6FLPev7WeL4sTFrqDkHQ8
gToCHrOj6/qaMt8/TjM2QaEb5btjJE098GWoZQFaspljOdHXaeekGabR0XO+aencG6lqxQmXwOoH
cN3H5ZOE8JPoOtP0D8payfUsJG0mbqJyjPa5MnTMpOTyg9cYQUMyrFpM1CFnjA9pexueUDFPad3E
kzcI0CX6r+p6sVIWn/GXI4UkCHF8bMsDEoBxufJ6fltr5jdXq2ywEBULgi6jGEFoylKlfFn/ewt1
Jr5fLDEAwcehSEQ4XoqqNWif8m/+L1rIGvkk/ApCixDBaax4yo+EQTloWXDEw5yBv+PUBfctUILk
lrqW3VyQvDfFFVFs3PK1hAkjiJwNMPR6qaQqI+VQtInJ0MA1fGhdDBTcVLTckLfMcrEiCuJi2cSO
06lrdx2B9Nl/Pdlcn3ZQEGtNRCoJ1xKTuOGs6y7uIWP4/MuOG/yK6qnuvQD3FeSHFxuFwA5YW2G+
O1Ioy8jyHrpqgQgrZSyIKlHjc9CcNvA1fjQB2aSHMLqCg52r8jMCv4dR1EO8tVyAyfshV4lj5b58
aN5l86BmI9etjBCacKsObgM1AUpETRuPdYaGueBGIMW6lRTzSIAM/0DEOX6mQxI7Ict5HbVDfckH
0iWTnrEu7dpGxgo4tgOojb+zFmqAsVyLXWIKT8cRc1mM8GOppb3rHKbF207N65hA9Yhx7KGxaqwV
BdBIHkGMmRYkW4/AVUGG/RVuzTXeRuB1x4KO6tp8/aldqrjmEgYvZRbVenikswygoZ00I0mt8frb
BkY6CL2VwZNgeugnel83aMiVNM8SUuD/c6VDfYZB5qcgezoYaJMNnbgk7tSX9hbnRG5Xls4jVKMd
ZDKcNACnuoCxgd1ckny05Tsg78EnmANNvpSnHo6l3HUkjEdC5uZbfGzxBgvQjLbLqfAb9gkywX5I
f9HxHMBVqC9dhApXp0X/dUr8kWw1M7AhSmz7HYs1OutseFnDUBJJTvRHzgKBwTI/FbJIhbwHO3O7
M1aj94STGODvtCUVNH6xRaEl78Te0Wwv3d7dciRRMobo8cRSX9yUuwbN2mDMn7Tp/3rwRuZFaYRn
UtNgdS8Ldvn4uWhs56V2kK8lE/zCCJFFOPNr9loldh5Px586XM1Bs9Gm/4CrIhsEsUfsuJNfFuWM
T4Otg3/A9ihiF1Ay7H2UEgAopIVZV7hshekRd+POuNKpNqm6EYQ6NPAak+iYTWApF+Kk/TddRJxc
bwNawp7mHhWHvVbClMLmU97JSpddLFFClUa0WVfwrh5Qe8xDGF+YuT2qVnhCHKHrmQ0d8F2WSV5b
o4O0cr9rgQtxuzmdEco0R8448wWzCLMVQDLv8aG0V3JXnWvOLd2OCvwDNGvue5BonvUo5J9AQM2l
V7n4r0npxMBDa0Qf0IlXlnnNLzSYHn+2PhnP0fFU9rp+dBi/ccI8x5Mj+ee1Mec2kX7723OLWbaj
wj4uYQrzVKccTH41RLeHjr+qO81I8wf1+Xv2kXuA66KRUoUWX3qohfeOqf1ssSFcgAxsb1f3rxOy
5whk9hGGAatsTrDFZWdZbzr8QmB7KHVc+7aNoV2mZ8wLPmP2upr1ywHTSuAWhjJiCPpPCDql3mA6
N+Q6cRu1uaVyCK89ip3Ln5NyBd01nKLYq7fPA3ToRf8bN+soW64o2QqUDWXiInJS/YKDrsagw6nm
ysDgRq6yGQY5TWOg1ZXAC2GICX4azVN8boU4o0vJNV1PNKxQ4QRQGB7cNtH91DtutQeHAPMMgmmT
un8DgOys3+j4PAPeON1HS+rAaHv+xy9LP/Ga0eDBpMagUFQX2NSNj8Wb+2kEt6MgfpHArCeC9683
X91oBzaOvESsMBRpvE0r7YmRtznDUS/X/NUOB9tmqqRd8c+iVqYGaBfKIcEAIy7bSqDMpNqrvQVW
H4LKW/l59Yg+4GxtlMNiv5jtlxf/1C9FTmGEmlWoLLYWuBhbnWW/tBCsvRcSaTKP60dj4hz+xzXS
aBWp3i37AqyhH+Ea3UzzXPVNOwosSdgMqa+89IWE5NwvWOv3JMYqTLM3p7mkrhlndkPwmBVQ93/l
pEDCBXu1OjZYOVrO9rldsBoreLCgKixU2F4MEXgSngJGTCBnZg6eTyFd2A3v/fuazbwmm3fB28s+
TBH6/N2FMYhcSvYdRGNMX9BjxxDfBBMK05JrFFW7BNEk1xfSjNHwet51DNBPrvLX4qkpdnJxDJEN
SAvMMqeabdzT0UyPUQkfPOTW3DWukp3Bnv11yYhbfhJzAw7I5KcTPXHhjtQXdJ8aRVdz7w0h66p1
i0SybLztBZFYOtV22PYh+6JOyQuj1L2I6bpbEt9loXvNemvwFeI+eGbevUB6k6oPC5suqu0XD0jn
jWezXA5TXSHTL5RFmQf78YNLETq5lX9cF6FxZFtCWZqWXcZTSkAcuFzc59Ml1ZXqXXV/Inhv6sB8
h+KoQCok25znaZuN1wywCq3+mpRMoLK+pSV2GeJJWN17AfrJxveaFb7m3lk9w0xkYoRL9HSUR3/j
E8sFiZ3xQT34D/PgUdQrwPM+9h4zH+HRxDUMZAPdGmosx3y9P0BwW0eRUMqKGH6uMJI6g61RssHK
w1OQeQceKn64GhzH3w8bal9XDmo19JOGx5papSuJnIU+ZwXHtTVJctgDBwVmOyDV0rz/4DugLlsU
YRHrBRD7Gv9MgRNr3HNTz4uSWmm422nN1s3ZHXoaySjQldzdd7Aim6JLKpYujgAFA8GdhWJCw+LQ
bLTGp/UMA09z+c/pQAXMxDzDyVkkpZdW6JeNy1zi5HPEGrwx3jMjEaYs1yi3iiVtBMpycFDu8/8Z
c5Odz8CsJoS8I90s8UmFE1FRSgaFP0gkZsIu9lpfeD0ft89QW3aJ2l7LFb1QlFE6laoYbJBtBdSQ
XJyxMpuieT3xEQug3a8w4fPcNzXartXnXObt/1LraEYHFmg6nVCSk3ajhb7JDPGux2AWNE8iEa47
mc0FAuzUxNAtE5lrOlIO9j+f0l0B7y+NTwmwy6Uo/1qLMx0+PUkoLuHSPTUyD+/dZo2HpkHLiucp
LQhd59ObVXgJ+R4DnJBnbrg1Me3a2ofqeZVOoGzZj/KaLlQPCxgMivl0xOM5ZtSP46aXHo1kmSJs
kPynzJD3xghTllUPaYv0/uzc7/ZYKZzJj+fbbndbIm/RYPtAUivmYjktoxNPn6o7wtOfEY+kZm0h
+OkZUx9ACq7M1N33PnZmTQQFS3NV5jMkr60KpByzaF9g9oyB+6zd6vXh3q5mQ24xI3D/VR3mM05i
mSMIRuwgYcphUg36JBaxrnIiBRcKDYRJkOV4DF5d5Y9XS+Fh9hO12hrHYfaPdYcrStd+/+tmEIgn
7XkNqsZ9gYHE9dz3rcLNTJM/wyFepggt3Kn8tEXZmkvQeYnmYKKerHt0AXNaYLmdZGHvnugD7stI
hRG4rupZrLKcZ6rDJxm8HJA6gd2HqoPS7PRZtFr284VDLrGcVX4LHie2e6Mm5gB8YxYZI/5d4nn/
mF1dNRTEics650+JEuoqaFUkcX7cftj83KoVuKPP87Ylc9XOvFdjOaGs+idMuP9yZ4BxRThkbGl+
/v8SD2G25XRzUsWOF7ISFRP1UQsegmrt5kIrd1hz4FQ7WKSBQoSU5kHb0/WdyaehaRWJNniD+mci
sBXpEFru9rIdh1H0w1GFgy3aRl7PNgcJXyMWPuoNoSQqWynkHxnWooCJ18HnrrFhag29vIwcrHlH
sIaIsYK5DaTpPiabcqY2xlxPoq04B2VBmPSR7jWDjGEbp/PEsoTFzxVW2vhJrv5D7As+uFXTv5FC
kbo+XloG3DMYEUeKMh35d+BQ3iJQGzdyGn4iz0UiOz7XRCecPPzvAsYa5ts0SKCmJYhd8DlZY5jw
Od4KYxRyxYAM4eLJQecoxIv6Ip0NOn8B28X8RFqFdaq/xmpnQ3VxEl1EprKXZFlJ5aUDxSBsFAzA
t67W5M5gKZhKBYog4xZfTe6cp4aNGY6zyV0h+avhup/o7IfuyoZYNJ7VTALtm9NK58jRHauTOVmn
g4NsUgS0wex3Q6CXqQQ13Qlyd2bsgkqqANZ529Wc8+G5MCHgkuc/2ltXeVrepxWOAloUZRqS1wA8
vk9BJGDCOOz/QYxcRrj7LSEfICB2ZDYdveRafbMf53achdRKawKCzlTbjSF0w/Ujiu1lBvuJFFL3
REe50vXqU42i6XOxlkLK6XHbSrSCX8hiDcoD6W+GA8IhcvF7nN/W4SYdkWcbdu74CQuj4yO7AQYc
b5GBvGWNQVSz1J1iVSVI/AWFciGvSUQWcLv4dZWk6dFmFsCB+l4T2biuKjUW1b4IrzVlzRWOzRJw
co7na/c+ugEo4JQqC1e8/mCuSxbWL8UcLyiDwiUfaNu/fuaYVmHx1D4ivRdoM8B+3bDYfY3RNP6R
bWBHd09MhIs8XZ9DR6sg9fLaVaD6xYDEJ0fH37GDBqhykWZ7WG5Sv4ppru5zHgSAcHUp9N2AN71s
Yf0l95nyu1Poov6r6EU7F8CyzpMvXlKTzu3ZMOQT0DJBVqlbjalBNJGuoOY83gF7Oi2EW0q+OZB9
5VusAGaScxW9vimQui3k9yJ31MZUNXovKOp4tFrBKmhe2DAeBQCNP7rmd64vt2HlkfV6XkIQ9YjF
szQfUT9bP6omKxrsdY/h4wfnPC63dhrOLyy0YWetIwVAKy6dY+5vV2ZNQ5peVmq8lpkDItpoaJCf
E2rtGnG6aRxWm0ujRFEXN8vRVpmcEISIyuwjKcwunzlWgFphXW0v470fkGUMC26ff7obxYsqS541
HYHTMxXvWoa0GPzkHkWqzd7PhO0st1bMfM1cB4Melk7VLltoYZq0sw3qrAr1jJDeLuXfxtXNZePC
2ootB0qYS52cll9LdXyzFBi/f0t0Q4UYY0vFpUxK/HQkcf3bUN0C2QFtBUyBlwzvwZ6NbBPH78x/
A4aVrvs84XgE/dp0GnKqGFgqfx6mRGFNsB/3vgF1MSGRKtLQKiNMQldZ1M1hSY+Le091oIwYZGn0
cpaRifsWWCw/rb7Q0eW/2qtFSYG0BUsXAwkURDc7AkT30GVg8EiJvDnYc/oQ2W6k/8RNB1+KVInq
T3eiQpYgFe4I5ONS3Dn8xEACJ9M+oCpwi+4ByDB+fwyfu2ncX/aIjrcjPb0flpDuLsTFPbLIPRiA
9zfIZh5A3ueklNQJnZPS4mduZcRN3OBs306KP/q7INdpLydsE4LptP19jxeJqtnvcywWxyXmHZnA
YtbWoFN3VUj+X+TCDzwWJYrq8ar0GDAzb9THtZ3V6wIbLmNn5Hr70+CJjf/PZMOazo62cWrLN2MQ
/bRlGE/EaVpXNeEPGjwG3lMwTQAOsMMWh5qqHhjEQdhqlVd6zFevZ9oUP/6/rTUE0RUw7zLeqieK
XOy+5GY0bsSZDsH1PNtwRhk9WTCEv1O1kbVIxN1zpu0eaAgMDcJgVy8kH5jKaSoWctkmGkFPR1pF
BvxOIEZOOSes2n3rMRDB13cpkuFc17X87Eev8XEVyv9/hdjydyq4Vm0YvJohR2sZ1r81xM7k5uRe
1acJIRBHhq+9l6UQ26t++EZG6pyZl+E2jEZb482ZBAD3VK2KKj3qUA6qV49IZoOBu4ab1rcn1g/8
J0K+agH/5cXPss7PKYxm9Oq/iAXCeRnQlADHhythYLuJdxGJV3b8Gd/vXuIC9Fxo1u3rj4JAzgw+
qP44bBsBfhVNKa2YkY7gX/F9QS755i43/iGhGk7U8WXy8LB9ZB0hlVyO9pVpt2RX3CqUC+0lORUJ
/fYsPKxOs5sebVcR3FDbfRIwb3hXjNecvJe9WkgyKXMcYUAkWBAHNIhL1t+6GVXXxLNdXcf3F8Eh
vxII0ARLAUPSUIQ8RNhG3rfAIqqX3XQf63P46v5Tthi0SOTtwmyYEEDRKWTMxFBy5qayYJEkyxpm
uYEhJCXp7FM55KxAKqPRvFE1sIso1bb3DE1YfkONT0HFCh+FmJCLmSNWcSWRxmuj09xTcSmCzY3V
e3R9wh/P8SvfiKXX9mqgYxB0PJQj0mR6S+/u46cCKzu9+xjWAfr51AAQIjZhleCESMX1KolDE+L1
EE+NblnkgnFI2pu0chZ7RuyXb9eCw9UPjzJ2B6IXE4jIy1t6CmcFJPwrBKtFGsv3xThuWAb3uhls
iYNxOXTbWxvRyni8EMGE21k2XEVjWxLbrDc/v7ED9bZgCD6J0nZ7FGtMagcO09ACoBAI8CynfRDf
5mhGYC3xVgh45cS5OL3I2T4i+4jciDXDFCCHr2r5SNdq+CuEJOisHK2WO1qvuswV5zbm8PMiQKKc
xeieOIRW5Y7yvDWza9Ft0IU6QKtZeicH6HScl/nNpJFoPQfgBA0Vn9N5JZow7coRQ2NgNKsSxyX9
QphnJojnMvrPC1EDaXo5ykCgBLKsfDXYzEpLlwwZrncScpoGAS1o8xSQ71Rm6mo5fLN9Qk+46uAj
fCPO1ePk4RswJV4sdKKUy8Q+QVUFiQVrJaeJpvN0AqQYpN2ZyJ2OifhJXeWHRN4Kdp8ASoYvBfzq
OCccY8bHgnMdc8nCi1MrydNoNdARMCmvN+SDGyTaSRAk1Q58kX6+oGiNMKNfPldMOV4m4k4xTx2T
gPlFXI8zrZiUvpsDF4E+naK9djKLYaChgOcE6eQ8AzSDCrnUFOKJBwXm0ji+K8JL1rSu9T+osq9I
CBGFfd23J7kb48jN7lQIF/KGraUD2Wa2qryX7ykXthrc0bynFudwLJ0d+rLF7Ronl8XdnfEGRhtC
Abi/bYrtHS+3FFcCyr178Em4X0Wexb3s18U8iqWjXYoCpTllbAFzKoTrRX/ez5Wrp6sQVsUK9E3m
9TUnFhzUYtGzYA0M23FDo2/epIvdjNjI0HthSYv7lKm4bIxCUwBl+Kuij33+/kQHDXmzUwDDL8O3
fd7gus7yiISBWXo84ciYfx6UMk+qf5KpUYsHTwOdtDHQZDuV54G+9TWJATLJgdxXsjMtJ8nBYQJv
KW5ZCYMbg5CV5ZROE1u8UiugvpTP14IScp4eUeZePWUGgpWc0LhF0Ef/w8QjhdVTZSWfApt0mNsZ
7bmz1cpLEhqCGCGBzR64nYNrwPxff6rH4kJfYfV74/f643LCEM0K3IuP5DMal4fjx6eTMEELMD0G
SGzZi8AuEqcaydNMNVnqU8WGP9FcJTNEHTow/a6YUgBvaHp04jKtzTlwa88Rbr+kpa3NWfL3734A
/BV/YdlypP1/wG9C7e5AAAdxN1VkKxJeMG8D+k53Isv20xilJJqGXbE9qqlfKAstKOZS9G8tBG46
NUH+GQDEwJu2SE0hvG8xg4XyKHMHOjak2Mf4tgTTDV8n8Z6CBXmqwKTLqClHgPWSp4oXxjJFrp1q
UY8AjqhxHDnPE3dxDx3YL6HRmaKoaCWgWMcX2/b4buade0KeBOi66T3JVZxzZigaJcEijJggNuoN
51RstZHNVtcFWLaunC6yrKlO28Ps4UD9RU25kkuilmIb6zyB7E6NbSqROnge9OkyIzNSh1c1Qyyb
7GMdSQ5rBlvxMdMLx9WjkuvSkTfao1b3I6heWL5el/ZwXgClwf3D+YsN5XYUHkLaZfQf+mGHVskr
xOET7G1mNvxRpFtTgxDIAXPxI8nWFzKjuzhoKkqWUV0ylX1tEGeSOthN5emb8NcTdKhE2KgQYhBQ
4wnYrlo5zG4m9PZ3N1zdgVZh2ag1o9BPrN9u1oF0Sza5MMWk5rCSl3cQH5fF5ZGeXGUwbWV6plLO
k7lAnSm/XQ8NnzQFcug8LNf6Tn/2uuOW5i03QTmQ50/6w5ydBY3WbLsaL4YWUzqJGaFES5jkgvoT
oSZRV8l1n4ONhuFInJ4KRKnTVwOlLSUKWi8m/Ov7tSPUX3R2/PjxtxMLEmiYsJ3ey6bZaJaW6afw
QxC91T/2yIY2jpkd4ErIRe4ZNloTEHL9cU5AQz9Ih/BlZsS7OQy+mFovWodfAIbanCUMBM8T4BbT
ycw4GOtYZZSu/DE7nzexM/9wTwq/nCCUP2qeWF32LlRET5mwk1W0e+qzy0KA4hI3edZvD/LwVYPc
Bifcqg4t9l2xTflqI5SbqOrl/xW0h+CFSAC8aXUnxjUOUE8675h9dQvqbD8sQiglkYdGEbfonLIT
koPwz+AYhCxiLW6IeCuFTeLFs5FzMe0nbCMRdlfkINsNh85p+1vm5ewofnWuoM44hBa/JeavoMMP
v1d7W3NyQtLe7s/wYohQNIEMEToPFpQtfmTPysHrBLvxB/YaxH9NcfmVgBDOU26nqpcgcYiHg2j5
py90LhAHx9t530sCpWlWvdi49WNEGKeYyKA3s7WsuYr5VjcCKYIyykhxk+fAOs1U05YbKKKwuocF
K2gggDf6+FtSNdiy1b7BtvCk7/Ve/V9OeoFjIY9vS4DEjrHWxe1arWAcuk9YPC02NB3ntpukfWaN
yfPUKew/KJB22Ffq3TM9GpCgWdwrL/UBY22WQ6za//LE3eht8ITj7FOM98HVOdL5RpmfZFXSluhG
/EkP+JlK9Sjag1xeCXyUEXWybtzT6blyx/aSM4u3bIkh9lCKkW5nJ4JOQ0G/BBdZ9DnC93Jxp6zR
8/55VC6MFCwD/bBZDyZUb2LyviSbRhGm8HGAW76SycTfA38/Ps/czDRuzYcWP5RBefLigDUMQ+Te
8b5x4KgYCqu19XwX2J9mXiyhxSQ70sCHjEr+d8XiE/ATlTV3qmdZ8beNO538+vtQeNGYTlHVXaFl
f13oBHuEQufB20evrhvFgFEvCb7AZPHxc4IrkM7bqJSbjzf5Z7IaXyaQ9eWgZ65YwmHw0N0Ndhz7
dxBXG+Yq4K64Gp5glNkhDoJRscWrHnn1nT2OguO1NAbeiAThbAXdc21jOxqrRaVFWigaMhWj5zW2
gBU2cpmJGRtCbdpBg3ZY/5b/h3wQepoiqvt7iub5wXEH3uJx1z0uJsk9Ic/1KD10/wfFYiZVW3CQ
H4SShzf2s67pOhoh/0fjbFaG7MuT+wsTo6NUG6uAGaFf/beX+CnbujWeFRJuQb2UEqfHQwP/Vdpm
Fmnz62LTnpe5KvODSjrSr0061sdO/clWMCsHjH3w2o2mwjnAOWtbLVECgmjRu7oQTSjAJ7f1bMR2
ljazaqdcY3f+5lJ2dB/LZaz8PZ6FWUx4gH5Wq3LJxedSfkAjrj8wm6fCNhH9uaq/uCoNcqOyMwvg
99Pvwiy+jH2DOvvxGemhI5mDkzwoo2Sigfeg9Hu6MgF8Sy0AAtNYReW+pb4BNfmijEpXAMn/6DS6
R0IrtAwTZ6wWrQtn5RuXKdW3yowKaIRyS8kztEI5z88uSOQezAnv1Jmsj+q6wXPRSj/eoogdslmS
8vXcwM9XIPMz0kXAP8Y4U0mOjOsE9WMExsmc8rC7E/jSS92ZWPqbA6OQcPHinC0Z6S32U6HRX2kE
rlQ0SejzlGLYdzM3nohn6SX4Vg+bqTyhooCF6vqHd3f8L1Gt81BK6Tcq1GpdmQxcko6/wj8hKsJq
aQah2wbOae0V9HmUX4ALpQobxKY3lRteMdhavel/+kQNJzcGJ2Pf4cVQ9Z0lUHRMklvdW7e1/nIy
oYUm6rXdr2LkkAUBpptxcmGOQbRqtinHIHKZuGbdA5FohfyPHxydYO0wOZCBad6DT9KRpNRD0oBo
VvfNp0uyNr2aSHEftu7ZM39+0vjYO69xV76XZ6rQrmh+Lh5bAMEuituWMNfy+2vyL+Ci/5yQ8ECI
jhiaztYt4AbggAcBLHgNmADWnlZ+7vA+/NPnAqxcezRf/TnGRVjb9E+ZgF9oZSltP05OhV6llwDB
Ufjame932phxp4LIYbS66xXCMWrKnsD5gg4d0INKNu/C9sciXuaZ+Lj35I0E+Vf2Ft58zrWqdeG5
qvlqJC8+sBLsx854RD8M+lml1qEXYXHlZytIBYxd+4kjlvbcxj1xy7qpafSyc1ONaL8wfOUrzmti
RTJoYBtHXddyCG+R8y5GVs5pjkFx5iribvf61v06Z1ZoqAjIxT9zP0RCDWifOVARdb+egJZ7g6sW
sfqaB9HIPA6RG1XqJaUbWTnJ4BqM4+Bt7kMSicSP76Obs3P/fk6icpqdbbr2PQXpVpjM5CZd+1L3
gP4/D2bwYSoj6PK/m1XDqFH3VNcBWT2L3f0Xg5ASVxt9HBO9kB+vp8osuRDAFmR+1lUyIFGIvdod
x6dXYOH4ktFQEgvlraItXn7G/QVC9NqDetIu7IoVXTBjI9mGFlMSFd3g23V2FmiH87kw6Fw5qXaf
5RGVfSyBSuy9U7yGk3zOpDbUvIbHi0+hf10hr6B+tnawDpj83v/1ADWnyOiLt3encoOYcSmX3jch
OJ0txt5tLT7CMXwTgcRLXfBPrfHXp29lO5F2BHSGY8Chaf1rv1sK+IbxGvA1i/uPaM15qjzTXN5E
+YTrlSsawlpdfPOf0GjASSvCgj4DILkHW64OQS1jX49HWvscm5/tlXjHurO7YckGgDcAeIDAJBTD
o0v2ddG+EYuPwOMo7Yt5WL7UoiBZhXt5QK/PAcWcGTBG9JkuwcKRY9cmLCPwuVx2L5sLjHeCEXem
KQML9WD8eM6lT5t0mod4ZVVqbt/Wb7jbJUgtSylQKEJwvstV2T4T/YeHMu22tDaPD4MB/20JvPMb
f4M/vitUN7geYWLceM4HgBjmc7X5ES6yii+pUioRf1Vqtr8XOiPaCvq5ae8zzCTW6NlaSSRTesbr
M30K4UsupKfCP7qsw06mZDr42B76RdCkgv8n2b3s81FQ07s/oGl9iV7kK/m2JGpREs3R/eBZsKla
IsL6e8jcyMyYGvxHmP2y+H7BkY/t9RK8HJNRTvedGSeevFNbgEvrbNULKeCmjA8ofg2SGv84MCHV
MzEH/pG/XaRgoAdorYt2GOM7pWyWZzQo3vBd9vkrttFhnKs4/Jf2SobWIoO1xr521vRZF63eXudC
TRgBQrh+kGYtuo89KNMGtfkmWHQYF+30fAVRSBz4Snrrolib98gTRyFFpYbfddp1VenSWQ5IYm8a
cg255zKgeUf0w/wn94Cl4mIemA4MUnnrOLnCXodQbyMeKajy0J/WF6dMp3natwMfEZdx1qcGJlPV
MaLKf7ODjWf1uEIDi+9cVi71/EL99LfH2oJm3KOZ2lBk3Tg3DFm4GwN14DsL+nZhfJWt1Sy90G6U
hqWNQPzf/El9Mgp9XW0G37aou1WFS2Vdu/Z+EDbCyjZlZp2YKQcKTreKw+h3F5BMLM5ZMCH30CMC
4Sqrx2evQ+YQ5auvgKhFcaLXXSZ9X8xPFDv06Tj2kxFA9k8iBVRMXGe72mWR6yw4ycnhdm+KdmxW
SAV+cBnO/gSrxBUmisrWalgpKh2pCmwCT39BIvsXZuv4irnf+iArx5c7C69yz589449edBtA17Hd
4zUYwylYgiN4D0t0whCRYz4e2iqGzrL3HNhZJZG/kkkYKhdPb32td1UAtEuTkWSXEBXurf1R/Qew
PVgiCN8+NnMc9ZRUMgIU6mxDtGCs9KlwZtjG8prRCgqvR4NyTOwavVvSF/YZRJxfJWbySVerDIkn
+9/A6XqWiHCwOabuIOd0WdCLkFTQW5WDvn32h7JP7jT51pm5aHKh3fzv/SPXFJlIO8w4lq9+rWrP
H33UZC7GZC5nMTcHlghS4+dVe9ZisYzuxLZVeNAWYfpa9AnKmAZAN+LMKLMfF7LUksoK3fAYqFPX
xFRN6+DaZmgPhLnvvqmRkiPrn14i9wq/uZhyjd1szk+zM7BIE2q4sYkTSNJG7NxU9IBpM6KRY2Za
yxc0MQ4ezV0t/092WLFJFbNkze+5ME7TAtxpGv1uzc804fUc6ykKlbU3uVU6fGvRtD5r8ozVCLuU
58Au6cSx5fJBRKjVykboxR5GaQSRi4UlMM3DVFPPMLFTkoJlB1aaZJbk5mmk6UaiImb8L8e4OZYc
7x4yDVu7pIUvhEGro5aKMM580OUuS4uUkrPUJ2kp+eeRFVbOCR6b+iorCOd4Zd5xWirdcoKp3XKj
4W+hELku8eMzhGAZqMuVjbQvXy+PaaUMQAEiqS3DMBYeteFBzCow4ZsXyzkkRkD39ZdIQQM3yltb
jDcEkdanB5q8OavqCJodT5SG7Y6p3mZn5vsc8TTaxFT/9OK+gQkccn5lGGopgldQTdg60aSEO6+i
vTtVQ0Gxu1oUh5Yyv4UgoHpWyaH4xTMQ4R1z3ZbFe64yaH8dLuVu4EXmNxO7XMPI+MhDdgBnFspb
JH4aJMonRFP8KsVtSTwSoeKJcF2uU7R+Djw+fe71t5ktby0bnP7HJeuZGuosyUZZrvi+9LY89jbq
xkEQXpHMpWrUc3TMmi4WrxYPU6WIkyohNg12U3KGrdtCnJL34SIx586nFG9P/UTY9O44K1k0Qbet
AqfmZToT7EE/iM4yABfY6cMkSmfqzkfccq+ScJviO95MzsQ5CGm20VRqyXLNzkXfcyKdYKZqxNvR
dftsL9aWQURvH/vmvSi4GX1BDp1YWRhP9eszHG1si6gUSUjo6a0ssnaEAnA8fwMkO9SxpP49P2AL
IjM5gkZz0HzpMqKf3eUKWiDpl6J1ikVxTHgA7QolRrweWjSg6yIjfi4KjX4D4Azw6EpysfCQRqNz
B1VMLidL8CpAR3fV05s+cIDDiCf4zFXR/ynKUdpB0t3MwqVgrGvf7vFcbSAPCWb/zCSTgqHbhi17
Xiku74dNh7QOjMNbV1Xx/pjgB0uVX+kjoycrHUlz7qccSM+L4kDVQPH0Va+DsSU8ENWKNazTYlkl
d0iO7mHrNs77U2SsUaZeoVO/C32Dl+E8CupEizHU5FGW/HSzYvZx1L4UHFGBC0ws4VA4s6jsG/R5
Ief7h2bPQF9jgp3tbJvf9LDC61rOEX8q5ARr+fh3dlRChNDoShjglp+c2A24UGctsriFljQ1l+oO
oYARsdvLmHSziHDCTk3PWkwB1koNBF2EBKf3x1wCj3gsAd1a4VtU9JuhrRjX1b0A/NYjgdxEuAN+
Xn2CJCawJoNgXwpbbnkTOg8hjzEj/E1q5n9GYDJidTk8OKKN1KQjIm49lIzE9Q1vj0HRmdmM+y9h
a/Em1RJk/Lt/nWAzxwKRqSIvQoUpFg0cYAGvPMPKAJ2nR9wArMEp1+sNmvHuqm0QvdQQ7eEBOaRF
YmxUShh6OXOImJwX260oQByDAzhvTTh7a/oZGDYstFEyFQgwRNlZ0HZa5dK/Q9iAh4fAN1QNpwwG
aHKxkmqkfkrvANqCY9TaTjYke2yDAz6+2sHJESFDtkWmg4fmjJWEFn7qGimuSF1zaPKpnjWIjAzx
8C+B55YyFzUTC4K4OcmcHVj1AGcS00TB57zlJFnsR8G9r7K67Js59SI+G5umDZ5kATiEeFgNKZ5I
EDsbf2jnUJQK61PPjUumYStidxhGFAS2JQGL+546VVQaTEirfQBpLUk5iGd0Qm4vEk99exgUkWCA
98nTDCYYrcNukH77S0JByor9dFYeUgbCg1cGbfhLCz0SvHqF8YZupu78YloDwPwDTpSkj85oMJ25
8AfmdYTGZBjnj7maYRcC4MXT8YuRap9JCFfQfcItPA3w2sgbMik8VSaZ300EWT4XwdIHJZ/caO30
N16BBKnkQ/VGu8/z3LbcNyXGdYfrF6WQLWL5mKGzn+Yc0allH0RYSBQPjZiV5nxBOqdq3D4O2pj6
ILOmgXIyBwunmr4e58J0mgRuAYrDmbHuqOqd+yzaOPZwtzhKWEcp1w+A7Hk5UJD93VtlXC5FDFCy
MT0oXbyo7HxLKaX7P3vZoJammRayuJ6kOA+CK1s7uKlfyk17Cses+zYz/t/ODTgjLEsbDcGQ73hC
mX5a2w4vhvKi7z39TzNEpeD6S7WVZZRVJHn/LnKxNy25viD1Cg/pfpf3ZQ/PuxaCTbRlbzNRT9Bm
nlpcgI7DugWapW/RAd+6gXhY2eq83AQfIRKSsrsN+NWJDVhfVV1V55B6iyutu+JinD7HkczGvqs3
5WJLbQNzK9lmWc0Ya3BRw/GccLs/3sbGeVYPWAxEIPOWUKPG1KzinqQngHGZIeu10lvcEVxHFFm6
/sLXBg4TBImfwvXFG3QhcXQvpmXg/hwkZ33AEcKlsxozcT4g/2EmlZDZtdkmv30g6PL0/nFXSpXo
7cDkrefbPwhODOpU0spGUtRksp79Tcif/EGZWWIp3cidQFpaSPbWrVzRQMIe3qBsVBTItXKw9iHj
jJRtAyGxQ0EGeNv0t6jOD7pTkvgJoj37kAO5GKQzuiRgscev2XkNTH/NGgB50mNEVuHhEw7s3evQ
+wtHh+MtSuVuwx3tYFfwADRjeYYAvMz6qdip7gtQI+ZZ1td6UDp40xwyi6WTC0jc74z8IxEFbHP2
Y+NM2CoxP7i6WZ+f6J9nyUC0RMYVMYQ1Ii+Aou9vOD34TDMm+41RxkjKYIgjNAyyoQg6JtP1QJUg
qgaFpQgZmt5homCGOsJmBGfZomm9nU7CAl1bdF+FUNas1ODS5BXL3hxVBX3y9m915xCTcCTeuhAM
oQzODys/58AcTi3Oxhuet3O+9ZEia9DCzcN3hjsEguLG0NXHlnO+7rtHqz2Fmg4YdCe4A1D10a7M
O6ASUYKb68v0It2b+QY6hj1qauEv0K3ha9ipaqzrYBquDpbvtGL9efB29WC052fZjvDN7r9TOg9I
XWzO48izXLkVfOaNZ8p+CE7tGdTJol1Oe13Mrw58kZlKkQ3yRZrsScHXi95M9MOyayMrjJBVdkuQ
Gki4xdkerIpBMefGTouI7lFIgHvsfktiQPNWhLaCBXLwDoqoLeTasaNDCEutZTNRfPx7UKG2rUmE
lHAIVLc8BPa4in00S/jGCWkDLLRGMFLziEQV6H++gZbWOnc2OKe7vrPZ9+ciNVczFEk7zNRC3ALb
GLMdy3XtzmdJB8GgD62/5bfsOA19ZKRocn3EE3hYTe0LFLpVGAsW5PsBH/WWgUcNqnBoIX/1f8q3
W+WwxfU+zowG4euOQ8z3JEHAFpvC0risTlyFns4HCcHUX8vSOHjMKr4wWdeQmB/Dv808uwFnyMtq
cf10iAntk/1kRKC4nGufiOn1vyugF/ecMsc/jTGPWFKYniIjvfFI+DE4lfpDtbfB3quBa3JktRlg
ReGcla6gppQh1iGMLYbfN9BQySmMm0MujeMFAvlTil/zXAAL5S48G0rRymXc+8kCRdbPw961mRkV
3mSyGtx1HO3uhjcZu3XAcar1ShA/yv5tigMiuDOb/nDXYj3XpQblheLG2Nvi2dKAJZuSs5QOyk/Q
9nOtIJ9L7nwCycO2aYT7pWAmiaX/5A6VUY+sbggjV34Uf/MHvpRBcZOx/KDl2aFhqlhRFzoIPBv8
C/ZSE8+RjwCJIM6h29wNn4D3aOZ5RH20X+F3VlcrmqpHr3UW2GtoruEvPOAE0yBVs9VkYMmo3tCG
ujbenKK32Qr6orWpeT4PvUv1BDkvnq7Ck0tdPlUAKa2ouPbtDzesACBjY/1jRNy82K8nx8heqP8H
c4E1Gay3xGs81+eimYKsFBSpJRxv0Avb3bPZQ68v/pnEFXjjG2g9Pw8/0N3XePwJXgNpvgmb6p6Z
TNrgwSW9azfAEClr5zaZ3eo0A+QsONQlJSguy0yruJibNNdmhOIc1X2gXkP3IoNGmmGj2R5gMTnN
QhXuVbSUqLvWzmEHIXvJGWVSOgoHRt+FjgoWnluFXBSHXWtSp0lAZykzsgbiqOT8a7jFV2/pUTeW
lNwCoXM3reDMx0GG2S99O6y4rKWPcTILxJe/Btbz0rfAr4DfetxTlctNg7Iox8XIWozKdiC1QlkC
0LLkr1au9pXC0nxzaHZzIIPTZZQJbqUufGAG31kjgBTKO/k7l44PjrHiCwlC3WDMtlbLD09NL5mX
EiTgL49IexZO6WpgVxzasF5qwGJnnZx5Vm0jLQf06264S8gMDhLG1SkVNcGreIJ0vN42rCeYkGzV
o1Z8AB2eQsBJu09ARKgxFHCJffQDP7ADwGc+tQi9zbLWTH8OHcBE3KJluhGwblazgaRwur1W6pCB
P+GMDSNoGW82QIm5aWcjNQ5+LLpLtP4HT7RsPZWnFxm921iWVxAkV8pMxbVAIHi9zX53j4lxrz+6
0z2dR3thlKjq5tN70kmyoRPDcgC18/lyoJ14rPmpuSVKzpMu57k3Dl88KOV5ebcn2eItF01r+gLC
pXHQ0HecScMw20w2x8vmcfYxdj37H/QIV2bKM6RAAapmIXQ3ciy3K/J0SuWOqkxtfDZrRif4MoTy
YML99mqYMQovmPklFVXhkYBp1OgFHUEr1s8ArQpqs9HcDxSt5sM9OzBNamKUUXK7x4ntgnWPClhp
FOiKaJWx7yKMz6ojP2A/MmTEIuB9Tyrt2zJUEIuQYVNV8uwLFd8WDcOEGr9B6/C9Jmqs0N21Ih3Y
byPqOJEXV73YxJyT2rLD6N3svpzzmJittiVPNcVHbycoHh4A9cliMdzYGZwCrceftch9wcHaqTUO
XSDOsvhhCWztYBfI3lhFxKV6qVr1BnstK2U3eL8z421oOXqqsiPZIczW4bKZDEnAVjr9DIAwUNZw
LBi9eJPOUVU6Dnnsv+By3mnMxWHgtmPWmfV8GDAgTS4Il9zDfLVn34B9G95y8MPmQl0iTD2ajMfS
fff/WjdHx4psn3srDC4pGQFUBHUr8OJ0A1JbBY0G3srHwmgsUlPB4zCkNfjFlYyVjhP92bSXCb6f
LcFOo1Igh3wHYKiQkT46Jo0M0iKwncq0KqFERxviVnv8aIHNtjpdKja4d9mTgm0gj/Q/ZKmok6+t
pMdj0mG0qZ0ZiGBW+Tj44ImtgwtdcJJNYy8THomMUBKGQQF9qV9ZF/ZZlORa5UmOwzIIBehzlX6X
UVafbXN5dDVKFLGS9abkWRUsJmUp93uIQTl7D+AQHwO2OdDSLaNcJMDNjwz/PnIwaXaYPUlnF3FO
zbSxjUXZpUVg3B7Vv7TPkkgD/nFeuGzCvrIK1FNLIR3yl5d4VdQPsXUV6WIWIK5TLn4oRjpNte2E
z4/Y8wlBM8ImbTTtu6xfAT1Zi8Jy6iUtbzsIrLUKlJ6+Nppmf2qCy/h/j/nZY17ktud49IJ/yy9W
pRrJyf+hWufFeAfU9J791/jwD4r2y1002op9V6T4H65erUsW3zGOBH1fAdKabV7QTjr+0Od1p9j6
RPVbCIld4cs22/KF6FZ/ZevQCCbScF84wNSi1Y3jX/Ea2LgBYTyZEZg9nmQF7UatK77z+CjgnFQh
qfbb738FC6TwqQCZDrxrT33r/a65Da197eYvKV9cl9DFId6HmxOsijL7F+cWOwxP/FUnHd/v+sB4
moqNgKJWgir7StseOetP8k7OA36uxVc2G1rUarCxOxLNt/90hnpYktHe8y7h93xAupGxMKzEjs1V
rHvURGfYT2524Y9Mrw0CRj2vLbdnUpO6SkARQ98y0pz2lqcfxNym8h+XmYbms7C2iCQDEaat3EOK
LvfLUDDiM22hABNnObe3wc7/drEYW/8jg4RxFuQmLogCGL7gBx1G+zGRdl9ULnJAVJSiwAb207TC
sUeGX3fZ3W1F1pYavU0SpNtuj7UVosjVnofCqDmXLJeN2oSj0UGoXNwXFuZLdwQElCgqKLGdv8GV
1tM1EpQjr+QGNCr2ViDDtgv+Mq8eCXJz5Vjak3il/+2ZoTSBfD2UN5C37cg79Z5aMQMB6JZ+CDqv
SVu8c3x7L7hbl2H616izX61SnbwmqtSOC8xz/ule55pDoaYl9CH0YNVfboVTTrO0ycXg1kMnG5Wh
jjta7ZkuBqiNH0IAyHSJPikeaXD8lR2TLdxpeSWw5U8KSoubw6XtAx6GaQQf/pi7D7eIYF7ITVp1
9s7lBWAhEMCPu66h13KK3Da/Xz8jaYhVZVckD4ARv9F4/dLckGLZ24gAPdcF9xfBjfrcdEm/lHVe
P1n4ymrV2Qb2WZaF/qqMrQEeH+Sb3TiadxeWAWxic1S1rp8S1UCWbSF3wL6x89yp2gHZss7V8suk
aoYCYqel22lAgACZS2Uls5Lk1Getwol05NfhHKewAegAQrgWeWN4Gi8n6DqmK5uC7Djew+W4U/ys
UU5/qZ0OFoxhTEJ98wq3Z9gLk8H2YnMjkcpekl/4+fFqa3kvQQ6L+Ga7wBcovu5EuzdP8tNpVPzs
OscOz+PTsi/s7UdrjJXnS1m9gvI2BwOav3nvG/nRJH+xpoRjeRtycZz/YgbH1AcSpZ99o25Xh+f+
yx3QHk0v1BvaeZWxCa1UQgMnb3z0fbvvLX1rNBHSaKZRiixt8JA/9XltB2A9GXIaUf8PcLbNQ6gq
9D49xKRV86CV3Tim4mTWkQgu2N5P/p91j+xLeHyGy4wwOy5wCXLhYzbRSLajwV3NjWyPD60zdecF
4WFlznwe6tp0//mem7xEegRKVHhShKBHrb3FCv61RutcqGB+J9O5lhTAQLRv4sXFDyT+ZnhPw+22
kbgJcvX8AbtzB6HdqzOcU2OjBvZH/DKiZaAjumjz3gTMDoQn+2x4Hr6xiXplUhpUZeBj56BZtF9E
Vwy7ustGPHMjUVkea3z3b01FZoNzlSKiKwrYYZWlzxar8ZnMKoPxIqEnuqPxO7ZOEie8Um0rFksi
s81TRDMOgN1oM2tuM9Gm1Ad3137NssbUGZkfWkSKiGBzkorblzaNJSf/Y1wQybmfHxWxZg5DKvMW
1JW2T7GgNu+Ng7/XQ2n9fj5Spq5TYHmXH09U0XpGAme0aJNO3MCqJLiLocgar5EZn2mQA1yDiLLx
u6xB0j5ehtoY8+HtM0AyrQtVseru897WpuWMz6I4i6rxvs4LHshWKNnBpry3rdyai4lpH0C9FwR3
m5n/ZScanxp+J7/6dH8iubC9sKuwH04V/K6bXk68ql3kUpk9SIdCXUShrlDzCFGFdtf3ZCCS8faM
/wIde3QYl6pVaWpeeShK7n3e1ZRMna7y+03PBIIfTJ6khUaWYpdHKX1HcGAAPw9TrXhkP3pT8FBv
qDxzqP/LsoPCFY85wgvGBOLblD+C2DYzkZ4DdCtjVs4gs+cvvMnMW9PQdEjFtCSZ+WNO03LyJrk5
LMgrTdEB2z+J5pQ9objrGOj02fkF+hgDG+HxoUBVFc2uLTkqoOZxfIaqVL8izqmJ+WurqdXfjnbk
I60puxB+N90kByOc+PpHdCBrfvfW4e+Amb9XpUNI742qZfY6Ybn1GIAn8WfYoPwuRyKcCnfD4kJO
9hBfRa1H2XQ9QNWPIxidLj0fCCF4cLTlzQSwYAaj1Hca0zpBh/MfHASbmY/SWPORs/DngW3f+aEb
ZR9EMQaMHVZCQ6OrwHYr+1gP8gQ/l8S1rAMFvpoOTh6mr9iP9eiRZExuJUSrHhkAtVTMCQXKi5Ks
Cun7uciYMhSycfSTImwPs7v1Hk1HD6dVcgtKyHP+bURd5MGsxOUp9CxdtbFxMtrsveD60lJHxfEm
jtAxd4pJQPBkKcxmG4+LdJjxUOgHM7xnZf5nlTzm0notOgPAmXezSU2FueeWWJ6BjPfoCo2RYrvj
k1W70fUk8JYxBtdp9xC49+dLq3V3ctNQcpiotljDhzDW3PrrG7eajBKygy2NcUjv78f8dhawSQv1
xIpEJE7pgEnP+5WBidMpntKctzyT9mMZSyAk5HY6VyLzHut0M5V3lDwv2wOEK+mmduXKLvjHZm8E
wgYT19V1lnMj/5POeUUgDS9LJL1XaaRUEzNPjVRc7/H8P2zxb1O9D0yzchjEeyDPxPwY1HZldYoI
LvKoxwWm/eFgSpvM6UuTZvfhAqDUMQgvj+9dZrZg1wypeo7CzKupplIUE47AnCwCfAJBVKW+sFwN
nRO65vb2Bx3qbdU7iT9ePEdVbj0M0xGrk1S4GvIrd6eba0IYg2nJuWP2K1+sxYl2T8xLrasFNGRi
T2dP8E1IeO9y1h85TSqnWMj+/0B+DvL02oc3OK9Szg6DgfZbfS/SOsIT93WVU7TuziIHLHEiqD9C
RVZgJ2IvygovAi/gtAzf8ySIplmckKT1KbsaHk4OOTDUYA8L7A7U/wVX+kpMLDRl3dY7Hw1BakLK
7MG36NswGyG9xR/phu0/cLI8FJ3LLlgZGWI2D8A5dUXvPChFGh0aJspbANUMSgg8XZhYjXXelNjQ
UQO5xTJEOa1XTOuNpiWkXmMZlLsRXmd+iIjD6d467vlycCuGrqAOmIeFF8Rl/ToIEVseskS+BqtW
8y0GodhNxRbWXdweCoBFmOS2bTXBTq9YzPJ9UyOHevJBXZs9cqUfgbpEaB3T57jPKhVukboixaFI
Yl4RcEoiI5CGt3XOnoWdZb53h3bcDKypHpmYwKKXbngp/EHQluUPF3sDtfCz3koClGvIK2ekcGxK
1Vrvm3eMdRhMnHUzXjygy77AwxMfXuXZ/oDU9U51ngRuQqIvlockC3GksPDrEVlFXailJgVkoeCY
le688gsZFP7Wv7Dd+mXg7c7phKNJGIPOR99Nwj7+Ui5hJ59mEXj05wSYK5QVCu+orR3F9rbODrFT
lSYnLMJPRmzKbUXez1TP4VDQx/jdAH+rCY9OSjr6m+QhP6LRTKQ9cUGArU5Ba4VG/mCsi2ePnYY1
tGPXXBeVhahIzm9CjNmRapIMwVCRLn8/aLF9K1g9vxT8LJsAJwvrsBmPOvTa7GrxdF86EdohV6P9
tMD2v3ekUzTp1yasBxP9LoL5paSvvxxCeZHtI7y8IAg9RAXHrzBA5BU17cQUJNdpfzow5yt8Yd3J
mcmuR5JLvjtzQMZr9MdSZ1ycMz4RR7vbk8GKD1uT7W/mTX0iuLa13f8+agZRfUUIzHE+fV7jitQt
st1OP6ei+BGs4tof3WxdftE39P+Zb/k85Poj+66PqpG8qmKHHCax5kZW3ynGLqKSgQEtY7gzept5
ny9cJ6CbAyUQJZeMIrc66QfcH2xDUiDn0w1ZszCfFZ3jrG43IrebG/04G9dkJYE8+QM873kH+sMc
1uCOAnBZ0PAWxWoweOQx+lQAZdjUOIfU4KLmMrO01Ga2pmE7TXsGN4vTA68MA/j77HaODvwuwhRU
44W3z0kSJYBlS6GikYIzXG8zhyYCR144VU/4V2ZzC+JG575kW3PjNo0LBlu8cihIQ81selIfkjWY
oVizPKmZBjMvj+022j6RuFhuiQPqLSPeV8RwAZGRYRaN7chm0aCeTg/cjxUKNNQTFU0GrnGFTgso
Zr/OukV1/4RBZsFTTf8s4edtqXQ2WyOFgCZbC1ORpCKavRxjoB6wXmREN91jAb4tP4QjlFJ1pPSe
gJodk9piPJM6ezf3TYMJQIpwFrNvVbNfKcs+oglk0wdylVR5HJWJqOB8myo9pXe0/E0sFixTjfRz
Fq094EKvcI3Gtgidminx2tpJMzC0Jx9lJvi8MaysDcaFg0dFEBDgZvSNzA3o3rpbO6l4SOzRn7SO
qt7OkgkwGDPbovMoK6oq29yA4QqQq3yojSohhMczFKQWH2Fogpg6wsMEBHddtqiIdOdtjJk1CDgj
bA7727lN7WRFOZ3o9LYILuc3WaHOfrvk41LDjC2au8VPIMn9Q6mprsSzSa5s9BkrWdq0WgEtayTh
02OsLMJ/U+pUcGX+bqd9lPPHx5BSWQgvgNyxJD1hu8SO94YeClvWOANGcMSyD02qG2KAD7V2vLlX
+vM6oUDOw9sXROcYzr7KlCjDWIHQxZTYaD2MCC45aLjMdVD9D9Ormg5wU4gxClEx2yYzxCJUkS3C
89J9A8GqV7R/xNtY/XYTj7QXItQT5InDEiGptZBpocNtKu3fcXLrboAojL78mLh+ic/L0fUPQb0P
uYjIfn9SyoOsnJuJlni+K1z8C8HivC8ftFf5iWjuXmWMudJ0cYZEL5yDTZ5VZOCBRGDUfyhol0gK
nUtZ6O98b3DMZ/9as3L0wxHWlGkz2DSSNg5jbe6pWorEajWobZIvcRNOef+EfNozyHgc+4d54XLC
82ftzUu5Dp+fk2PZSoQupeOkhhqVYcv1txnKWjTFimBTjBZgGoPaUzEFgqmP3NIrh9225U/f4nxC
n0NNFBDsJEtkFG28xuB3YcIkl7Jr/8dgaBoBwQHCzZ6TGaCQYduD1V68qPH0qNYhxDElD8QHpNkJ
TZyRaSrqf64U8x5Uw7/ivoDRqitZSYISCwKrQIL19G4t/FdduY5MyvuNeIS53aZ4QUqs3KhQlthu
uHLfTLO0I7uzeefKfa07rVK8tgqllVPt68FSLThK06iqSaBbqczEWZ8O0dYiVR7NDwOnK0kDjukS
n54ZMSzGOogg4j4sOFK1g0RlUkTIwziN0x85haryXsDGJ459GI1ngdTWvrejTakhor+pG4mugzCo
OxMsabvWW5mIYFl4pA+seJd4ViW97XLRwuNnbLHKvblZcmlcl2hJ5FTLQ+f83P5i4S4nL9ONn0UC
LRlPXEREyP3QWya3+OhgKPt6n/pouOzh31e+3GyWWv8Srfdldlz5c29qb2icW5B06a+gm6nsAvh5
JfpH+9dChII+Mg/pzGjJUSbwf+OT/aWTXtubwHM/Z2cC3R90iow6ETwN91VFB0wdZIRkADI+jK3n
1ihltSIGSFuwnK6FLQHvG3v1EpIKnnxYhmP8VTOvveG4VFDwr8ToUi/WI2Bg1/54L6Q6ocDNGcP8
fAwPfUZBsYxtVDxXXbD5WhVz/wN4pXQZR6PqP9ZP1BXNAVinm4y8HPyU4mG3aVjg93qfP5mZEwCW
VXSwpWieJ7GEmQKDV9Qi/WKU9hp95Nq8jnkY38Sv3ddh97i5djH0oRAqtYqjT9MBKu+NFVzVq7Yn
jf0g/OxcOeZXbmWYOdL3H6XQunp1FNVGAJiXRMDtF9BtNIOGxti8+UooPc9sKZwPFDx1joTsBu7z
rt6GXE6ak0Og4pPFVx3Ckg0ygYl8Vxj4ZaOH7TnNdd5STqfnt9rDud+qD6wvx5civb9e/h/Xb5sk
8ko0UJYegkmv+9WKIcj9PzqNkMD6ypGnhS9m36rCg/wSbxqKGj8ZEeVu9DM7F38jMUf0uQ94Wimb
wqFDWOmuMjr3MQvSvwHCNZo7d383tE5j4oZFnlf4g0mSU38WGQ3na7l9RXfFYJvgbr/JQpl5at3s
7k/gaoLRwMrPsU8IZT9UUdOp+ft2YNjmCuUVHZW3ZwJSVuc/ZB1UYPcov7If/ekpGbMnTFoDdoIT
wSU+ZWrmwsMEw+Ab7bD44FdNVbTPvynTAnUoSkrZYDcWXxL40qGer4rVDG+CduOT0cAwzY7F5J/w
RjxvebrVFVmvnEe7pcBAqi/yHo702nNx6UnJjFimxWmlnWq4x/yU7bGSJz+rC3+rDB66OTJ2kRsU
FF91+I4c+ZqLeqprlf7wUe/mdUQG954SoYBiZLamGYfQ3l18ZaSigsKiUti1luc0QEApC+7SsVHu
7kF8fAZfXZsVYPi284/A9AbPy9IX9q4MbqttATA7aWIlRxVceJiV9PyJg5cfR0kNUO1PV6smI/Lj
Lil5LAtH2tijZmGLlKdygr+Omnb/kiY4sVfDuvq/XkCW2pueoW9dnl4+c92jHnDnTIaYY9XdcGri
Ayh8pykHcWZj9cuJGukiFd7cvoCeNLVdIBXScQf2J7G7qS9RJLVYATHVzIOSOjnKeVJbSNKM5cIo
hJRbc9qrRhju39PmJJPBeKPuYsUbujjXEPszVVGRZQdTjLDDCMsdklvTXrCuWbWfMjSLqEe1cZWj
h22lSX00tCjQ/FZjCL65ctVgMAi2Dkkd+yyOSytjAhkfJt/Rf4TvKLSho/JRLMRncNtCrOkGkdb1
EuKdJEZZjnivRVijRQkv21OLQsk2n5jMaZAQlB8V7K0dyjDcKYDvsVgkHDrq4TOz3GobaOb9hgNe
Jai+x67fUKPJTf+ZKu90gT0YArVqSAAZ+EQl2O89uIsQwVkXj6KdAxLxTzhhSBDCSCL9WmM2mGAd
OQWqceWtWqkOaEjS4nPDwhmV1gsnrG2FvThqjrlONLx3hvSCT/w1horMeneOAZZdfwM0HDu5nCA5
N0FwjJjNye0U//lH6H6lxDrvnTkJU9+I59CKdmAiNIJW7OHNjw6eT6P5ExUKnXbHKI45wgX/IAja
wWVylH+yPvmeFOteSA7tHKasqTiay9MfPG8eXk5gNkI5yabMnPj4ChiRbR8yf9jnmznbW74kuRnI
eG1CaCwUrXnVAXwCsJFkVs+aLYvW7lhOjQAgVINHjMCPKBjhxdzG83jZhBdkXl0MOPYdgU0RVhsw
aM2cyQa1O3GOfjLz0jzvThzPWG6URaEdvrxh/2hHL7bGRfDMMTyAgvj4Wkz/XYToOoBq6ukkZ9uT
NQBpQ8GYczohQ/02rF+VFQSGxRkLhXoHOLe5KVAT9fWcLGjBe/Zqep0IdUeIxEPqUzWgyiUus4Nw
20gREwc5/vOeQxY/djWURDlyGnxppaYkYFe3hbZT3kk7TDvOZkr3ZF6w0SPfLNmyL9pGwytdEeEh
FeGB8a/Hdz9ZtkgkDh7YGt6csZNmoJdJeNOsO8Z6TcFzow9HE+668G4KXCbBfc6TBnLuNSFsmFl/
Y+2EQL1v1F3Ma/++YOrtuj/kjuKLonToZM7V3/e+3qUrmC8vgSUpAsjfG15SnSl1CjJbyG3Yfb76
dHkx8aEg7zSnk72WiiEqFevB9xlKSrdb3XetnlC4cROG2BKhTrfvmJptiPKsr1r/4/6Pnp2FPNRd
acJIewiUlNKAIxPrvITLX3EyLgdFC+uxqC2MScSLTWKUYNA8N/BOmts7TSHKANbrtLJq/FtifYTX
wZUdZJw/wqZsvyGFcLvcmWcxGiAk6fuqEmmutWEiyFOoRDeFf7IKZ9/HLF1CmIIsB47v+KjGlHx9
f0SCLEtWy7T9VNOt/L51ZgfdCEF+Xmjy6LDBSAfC5aStbSpc52RYN4XCtGbziPXsbs7LFAn3e0/C
yZ5IlNzzxKzrpRu3vt0Obzjtv12V+RE+VLZdEAVq+wsP+qPUcLjvupoqCpB6TMFPArjT0FSjFRKe
ave3FIieYqanhvZUWoRrO71ObV9YHDlRw6vkXeQZe36vmXfKnAsq4aBpn4wLnt6GUV6FFQMEFopn
H4hYZbbZ4rUfAQ5gM3ddeGHniwK5WsHT3CwqHRiwHvBwLjNon3YMSg1PoV73jxUYYEpCjnXZq7xL
TzBJYrRBRQSa4zGrrFji9JYOjyupPykO5JIhDUescbV/6WUV/T39yqcH9OcW8tygbncJv1RSOLxM
vPoyYKbB5g78Mb1G+qViJDMT1ceH2vP3Udkws0Avx1UejVGSh23vvVZTllEdSR/HoeAWdPWAd0zT
Ho6zVKviXtldSEtS0QoLkzVsPHNd10cS2Fo68PbSropWoRAgUI4PL9SrbdXylb4vUH/8ejcHBrUJ
eJ3O86ALZpZnHXpiInJiiiokikcTuu2g03l8XuH22yEGH6YbuojdeLUo6y8cNkmL4wVpYTOH+ODM
c8ssww9D/QZlLJ6ygx/78ljFl4FOkiXR0ZkAgS+nPuduT51BUA17sYbKK9wxkl0wGRIPUnsQAAUz
AvWg6802311eRgQqjknX0dS4/QZkGa7o/XIhrui8Fj1WL28jtHkF9ru28B/bl+BhhhU0ScgPRxIY
NpokKOnUDFdJHqrym1jRNlxrcvxhGgZQOypqpD/fJNJLlkjy5/it08fkkyWaEgaRqrFto465qixs
tcgBN8109eEMusfjAKsNRXnggSlYmQx5/BdviIO8OIek86GQzgDY1DlhiOqfz2uZng0CkavpjjP5
XC4t5n73E9ozornjtDg3F7SmmYdbObf7MMBlWw2k3Y7ysB4cF8Qf49WvRJ/CC6IeWXJdtkMobEK9
4GIOUu4HElKCriZ2YXNNZOMjpDZMNEDAHqJe5LvCN55E3q9lRYPoq76YtQbnIrWgPpLvzk/twx7a
/SsRoZLvC+o65Dvxll6mkQIYAcp+YX7hVmXzhP1f2QNazGFUpiT7AjlbNXM46AJUPJHz32UbXTxG
nuQve5QemQDnqWuDk3d9FY7Z8v6P+2WPaVXzq1RJ4x29rKzvfe/pbI0Ruv8gcMOnx88rihqJrQML
r+WNIHWwxx0ahHXP8TWj8I4NmMj4jem53dUrSpw5Pn6JTH6cQTVmkFRiazkHgnpVxlDU+pUqnm3F
Au9QgK7VxVIT5NVW8+W4YjtiCnvtGr3y+Ws8ZdcrMnQJAN+jFvDIQIDOE/c9sQP3ux/K7gFyqMLJ
WGfV83x9hAdHhJGiJsNokBoQUY8iXuHTujqKgccCvivts0liBBuJ9+K7O5oWqY1w+ScE4nv7djDG
XH4eZ/NlxkjkxwPq4PECpH5u8xEgyUPPq74xuFNHoxBwMra/cqfdGDQ17FwUGe7q9COPR/YUMCET
ThC+m78JbnhR85iEhTpgxayB0yLUz2coB2GGZrZX1q59kfV6wLALMB9CbkNtojah476411ohRBD2
azo+g2K8F1rAeKir5ZLllY/+vxzOTk6i8H6pCmhBQQAgZPjQSiikAUpam0r42JCqJADOWVoAMlWa
xopTh1uojbF/CxfGnePHp3uNJOO5qXCv3BbP2ZJ5Ah+bQzXLFE30EKDE3XNYMfONMfRufKaC1rXF
IgzqvdtFalZj535iiKrbG/1cPZ/IIvTBPeF0NgNyfUlMpTDSDQycWqTn1AI/ddrKEUnkB8s8PrFL
EzAMMogZ24CrRxNjtqGU37AkB5mHpWfKW4W59Aaa3WSd/pppiDRKS/8xyrgnNkdNJKq39pV2+Ixu
ghE/eyfoSrfMP5FB1vskw9mfaWX4TlL52S2Iu0I7Psj/oBbRiKAWDOcqdcjUsOfRkPKlR4XvfpYe
lzXR7aAvWcaB1Ef3JlF9ES2Z8rpFGAD0/tAjGcTZyu/TrYwXR60z+2pOqunDFWOuYIKpAxHHD5bN
HfSl/Jbsl40TvqHML4P6peTlJRUkrBQXhHIKqB/yq/1FoKLKD7e7qcUz30Ym2nTDlQNSM65CiA0C
FH9U2ysWH8wKD1qrNOOuWXZqxrG48P2CBiTbP/e5K45zgi/8j0eU4D1kuv1jpARMe9jzpQvN7/OM
EQ/btK6tMmltqK8ByuK+cDQnCwP4R1JZlLfre46ii6+uLJbG8D5fjUdEDCGhhAzpFAc5ZjCL2awj
8G2ZtF/mvV/+BNqHM8xGnB6NN8afVRNHhiBWSE0iC9p8HSKsxmJ2R3z8RX1UFrBJsM47C9dEDtKz
tZQEnPYFGNlG8qYODrgqibU6MPX8z4+WMWA5sscbUQ+4baYvWYc7O5naijAEOo7VfqDDayxjXQjy
5HW73VR4ERZyQm3QrKD7ogaMMw1qMUltGNaZG5sPPgyO5kJPTBGUbMzratExVN6ZGMgj4ovxUBkO
ojrOL1BGltetGqJz2tWg6AzJhiZpKeBcSj0TOSR0wUnQCPGr3V2Ppx2DXmu/HLTz855KGRRf135F
rlR4T6rPlvnN8AGrIf7+d2Ao9k414RIurynq/7PZtAfeVwgxy33JaogwAKwPwYT7PyIpbpllK4B+
aSSxIvRHf0I4Amu59+coW0yNbDxzbOnoSZTFUTvqSV26rtR+D706Yvib3Rxg8T9KzBiWMBJvTMU7
RjppY1o+KjuUJMz6XretjaYBXdNtyT3LM/cI/ggua3n8JUXEjWBQ/NWzA+e1ve+4i29dJbpM21BV
5UKt7A+I+f4dtGs81y0h6q4wVpym4bKLnUX1leXC7y4B8yYveP/ZE5ZWGl1GjytEYJ2+CcAY36wt
IQwSof9a8+v2yqh89xwnAwg8Cu2zJz/zYCQ55XWnbpGPq0SjNUq4IWKoVwJKDKvkSHv9lSjrplgq
GRr4el8p6JQY/BkORVoFe3h2E1uEfS+NcP6HuLn3BogrnaZfWencgOevzUR7dc9QhKFQENOtMuFg
eJR1bf8RwvS+QXC0MpluqjsaYDVeV0EbsC/mlbfv5cokiemBXCgx2aayejdC7GzInsAXjjcwWpYV
VQIIEcbd2gNfdqg7BwBuqYZMtTH90cgqbZTqz6umAit29LUlMNRZKfoWSlJAKJGQot8SGpLmMc6z
AHZFcUcmutaCV+x0PqIQ1V26XEs/fkHeHFL22wjf4dxfRmFNNZJ9NA4rrG3eHK4p7qQ5Smdc+4Bm
bzBMHQ4jrM25VKArlA7k7wySgjkoyxQszZ7Y++3An8IkaCSmNay51ccZMPjid69xOCRDGvzWKr+z
/mjniq5Z+yLYTsBxb0p6XwGwb+IILSotPfOlpuRnhc17pwWYvWchTIKN/1rAapMPe5kYl+Cw6zdK
LfvJm4bSWQwno2743DU6GwFL9xtXO4eXvJp2KCZcoLZhjN2YvHy0Trs/6epfZEbaOX6zT/OW19+Z
+ijuNLUjyVd6kTGRiMuXCr3HcDR4yNQYnRITy6gP4UV9LCUezMjc61wRm3zJIqhq/kszyysdaY0/
XLtXCv6zBkxUkPIBF6M3i9CSfkXy4XmnaGSeVUHQKBZomN2We6BAQmZc8PrHsx8LjRf7w1uIMy8x
/eRd44vO+cpH8KVlI2hG3uGoeucvOSJLGoFtigAyQYMMN1ajujxZMb2R9fiv2ldMlvU7VAR87CYc
U/egkESIc9ZVo6PfPH8WCDGzbjIJTLTfDcZyF6qI8ge1KCq/IoV4M9pEWhQaUAo5nw+bSw/g3kex
UTvzHM0E2kk4/O3UDp612hH5Wt6QqYrOr4m+Q9oakVi824e+bLu2MHovR3l3FX0PFChQ4LQFhFfI
y5553D6v9lo/+eKxPGg7FoRWB0yBLAliV4qArd5JwpUb0c331srYvBVi62WGshM6UmTpf0x+Npx/
3BVHsIOCxLXi7OxXL4QtwqHNrL32VFhutGi4xqgTmFidtxLfQK7qsHkLIMsbmwYRFvTyqvcl9BJb
nN9+Fwuvt7SHLSPZg0pKqikTblFn/tM0tDam418bUbg2BXlw34kkgwHB2CsV+QkS79/A+TUWHgM6
q25SaPQWFSNmZwZFhtYZASUQ2dxooKNppKz2IUz2GWh2O3q3ji3mwYg18uvGf0tMoE3qRe0cXzOO
/6MAtwPlJTNabySljQbqtRWofBzpBjQ1VvCFZdMKaoHrHmeCOLqWb8mZnKsB3KTAJ17Ef5Km/+Qc
AZcWADngji6cXuPXQCZNpKzCSzgoL1H0cmCWtTZttMX0Bwo14D5EQzAmbAnFq+Yn+L67a7/3chIX
whDWdmKkEkZhL7J/jCPS6eM5XHHApnz/qndeTjvEIwMi+SmX+roOu6CoDO12A9b+XB0rqFrFA9uw
kBXN3si7kMFdQbctPszSPElUJKAVkZFNuLZXBFYhmI+oIJyc4rUZ1HE6St6npi91gN/26t2exeap
mPf3rRt3Z0zvXVktTppIODtOMXZ9ycb0GCTXLDEFuCnjvrqMZn4gnAlYnKfP4RNkUocSfxjyzqhG
AFuulJw1W5DxZ2JssoAG3QoBWI2/tGgodxyt24mXQCzypgX2fRDX9mhkCQtA8B9iHFCkjO00X/DV
mcZQkbHXkzZm7fbJTKfQzMmwsDOtXn1Y+ecgpZrHNNoMdKCmLt2OuMZgGJZyOx0c/aUT6SFVVcUm
OhRrEz/0imDyGIiCjYjEMuc8Sk+figAWh43aI6zCJiCDh41r45QJrO/cto7TGfBr7n2tOPR9Nh2M
x6D7U+vPDHEqb5rCj+0CEo075bG1mmzDe1XgFohTfkdgG2HoWinlq+MM3KFWNOGhE3/i5DpqlvVe
Nj1I09DzOldvpswKprtYzDJn4mjvbeSJaET6QtL7t2wP5rNzgjYtYmsr5u5Ic68V50wOGSrkLWW8
xumDiNpYQWXbBwI1e408JIF/iRsY1FOnZ9JFMs6Av9R9pJcu9uFjQoZiC8LfzkR0B4pkLE3af2dw
aRYZqZOCzUdmxf/KVB2eEoTHkOGlgeNHK4648/kpO/PNI8hr3xkDOhaG/FqTJOZgT/l18ajh5h68
DuXrpmwmGqn3CALfyqdUEDcVq8cUxPzBDaNoLB9WnYvcDghIQTsuVKTkVP32Sc0l9RzqNJwsYgfW
FTPQRg1y5m2Gme0EhKWbWDlYkry9VyxvLnWV8UVCfUVP/PZkjjK0zswYfDt2QNL7z1K1RB3mF4tk
sdGoBuoUJvJcCTIuTAG3y4qn2sGMz+WEi8pHW73Q6staqOHprN2oLCjIdTUFFiDQxoVK/nqcyKW9
m2Xc9fEzsO5hUEV1J5IOES4SZR3iHXnq36n+JQK2l5+xTLO2SP77wpZqEcoIkHjDCxm8y8JA+JDs
+OugcTvFclomZ7dMiL2pPObd9hSWh8Y+ysA52GJv8w7OgO0KrYaUaiCMkQXzeCtv/xG8P24uvPHe
iXiGNEPK5hdPHnbBPpYDkWbf8RwODD4kR2CsVSGv2xak8cCmqkenjGNU+q19mSJZ5Q4+qx0NSckZ
HsvBuJUiFESYZSUgZFljvfk7CAYN24eQu7dwi+98ZdiU7ptfnOhIY96oojZhuEvWnsoogumvBfGs
PXDuK1zrqRDzEil7mfVhPijZzs5YuJNhktfTDDtBk5BFpwh43QVazuGnhblX0b0NAgS23dXf+Lp0
rFu/J3LpJSr04MF4pqZRe4ee4S0oV6b2liCHmRTwUvZFKeKM/bo823gt/t6PoxF+FPp8Th6nu4BK
EoZQVPnmuhapP+mOFb0y8+qAgWu8qBRkLzjpP4CD7+Wh8dSYxaBUGK2BovHZcp8qztXwLqy8S5rA
KXfT4aKqAd2vkmUHVpk4fxJDgvCnlDLgQxtAoxuEutWA6iHb/BwAkxwVNmXrgJ81ROuH+puDa/xe
7PcgbGHQvV2NPRQI2PMLU/Rbg7eLl0zNdT5EOyEsGi3ZeKkKqY9wH2P0NAA14M3CK1r0EYc53G0j
GYwfJGhNHlXdS4OkBzLRrXdRQgNlamaCdkAldlc3EI1oDjUkpL0slStG4x+uWVwyRgeFD+l+cGaK
S6h65dmgUU02cfYBA0hcG2bTDGcTgzb/N3HVmfDlKHGQC7RaR1eSgYypW5ytCUY/Sj3D9Ymqw5Hh
cVl9F7N7VJLwe6Ejx4eaUMhPJ/b79+9pM9xSgbgNgmuc3DcQsM5+Y8Co1Ih+WBcH0VXZp8rIkL+Q
5R3sNEYk7VbE2OfetqZgzzl6Oxv2/SB6yMT55j9Rr9azwPf+dxiFgTYz88T8/x52EJhbUKLLxWdP
7OLaXBT92tPw8B20FY9TDeHr7O6UWcRFEj7wGuHxPVwypsENwN2iUS8W7YjZL8D+fhiKUzyPZaiW
geLqG1au3QGSXo2NPdLJs+D86q1927jnSn89e16M/pim/euy46HhB+EOz7VqKSsHzK/gbKdZMeel
VuToamcCjcthDRFRPAOUhu9A4cIQ3BbixNNNjtB7LrW/E0JekOpbwa4OJPaN4dIZWOxzNAXFGbNe
WJsC1GTPY0WHbJLlmxpKYZqF8NXt9lYQqXpvFj/FNLiaf7QtmZoH99NOlciBQOsqdvJ3lFpq9uQF
Xp2qLqs3d2e/LGvv8sBMEhzq5xNV06GZaZB6f4v6nGTNbe8AwhisSdf4ymhAAzvZjcC5N3SwukjK
JxKDoHdk7B8VxtGGhBEtXJnco+oBO0yki6H2dBYnx7UlpGCarruM2eBTefB5IYN3OpqR8O6ua+M3
Wk3hJOjAsHa3coEr06WYVw8MZhpXbLVuZe7Kaz/nuTYrX0lgg8xyjP47eebW2dEPLs2i9CH3qNXq
aC7H1mf7oMTyHzXSNQBLXYS6KvCugmZlt4D5Hf+Bq/YO10hr+hJcBlb+PnrYAcIEgDwjewF0YCqZ
Y8rRBfgQ5JYO+ZncilBzPM0x9Sfmf/il6WYv1NjKnRYC2C61eXf/huQ3etJQEWrcZ70s05iF+87w
UmwPR3Sm/h+tHPOW7pDAc+xyKKxL++c6/zp6KSJipc9gMKpwB2G3g9jOGsi1z/tlL1O+IYyih8nX
sPGkHaSB6skIe/wwL7ZYP3+WBi6KBRYLlxyYfSooXoJHwFlTPF4hP4SF/mkfP6erWOtl+lOGiJNI
ckDburJoljinNwuESl7hRS7bVaKJcDtOY7mV7IGWC2EXJYPiAbC132wB4UXSwmOU1UfLC/yXN65R
MFsHrgv8xuMYjWuImk7ltrhKoHjTz146ssW9sgspyUMNGYCKfyByaBmIt5arxX6cPJ/tA6lubwJd
eIuyGogdLL+lvmAXWTf7x6jBklFPFnaaxCsH8IEzUu5bTanAjkJR3qVk2De/tnaQ9Dr4LznNMtA6
024uX+bc1L7mXWyu3WKkoG+vI3majg5I4IO+Xs7xcOUz5ld9l7mZTaSpOmgQ5T3ooKaN8QXA0Z/P
yeNKn8NV0qlpeGG4E1UkHLvJXuz9BJNvgORShywoYp52gpSABIsc4wNUvUvbII64Khst4f4rg3Bk
M9q2s4xQXsciWjw79rwY6yVGv1Q7Q667r/MTU4ASGc3oCKxGn76mTXYG8hoSGtgI4pByM5FrzW+x
vD+5pHWkpgWN/bOIPcOY8BR8nt6lSb12MhegqedeiVAI1xqajfQ9o/DIOszmy/MxKyc5iFWWZl96
hLrm8CSBsLDIcwaQvKIv3Axs7yEh5HATnBwpRNpuUFU4FYo/pl0+FNKjh4ZO+BjOOKz/JwTgn0lG
xdmtdQHoQ6mmrXrfR4ruAGX0NSFhTfyVdwPRLzKf+AX5NwDOUvfcixz9oISVb9/piV664FC1TRGR
FqAge0mjt3MNSDo8yyZAo+97+BQ2k/SQQ1RlARv13kfNdagBhSfmlwSUPjgMFEUOGWbk6CAhEhna
LweMXBMQTtmS5d61pyOXukJMuwUeiGzRpSLY3YL43jJqBsdment/O6j2Plw4luGQvzX5naEYpiKF
TZhqe9jhc/GUWgRF9Vqmvt4MZs0uiEH+QeJPYFgB5W0aTJOn7ch/rmuCVMFEhyMZDbf91Lhy3pdT
2ogKE7r3P4Ob/nprmLWGKyVC33+Nl2x5gf4D03kL5SfMYfdNocsQls9cfc7PgCk6Z+YV9toyWQwS
hDTIn6wdGKmU0RiAyjmW+1LlUVRKZsNJcEVDsANtUuSzbetng9z+Bo/lfIrtuVVLt9P0rUNRFG+4
7vMqhOA6P1jhti2PZF5jxcX4C3xIETLbWLcWrLxQas2JmkGOPoVrDxv5j2V+cjkOei5n2TTIGby+
SKpkSjtyp9z4vkcCpEK0owP+uCuHW6yQhWGBh3sAqN/NUNk4hqgPC6uBc2y8A5oqR1zb1VUzdq1f
sZL+dGeBrlW4wSF4oggTm1bMUcnM84zCFWssgYcGDYJZTMcsiCGVGW57jWo8TDuDFuDKcnmJEjxC
uKlzSRNTbeqIrqZYHhF0Iffqlx+FuCrkPBv2akNve7D6mqISfm18D8YaU1MQY5AjXV6PKfxHn/a4
O+06CT34CcIut8M9CVMZo59kCcRHxCq5jOOcb2WPM2qbrNfEdCqmEdTpwzGaSFMyHi/e6pVlcN+u
knK80VIVlb8ubFBubzLyMWjeE30T4bJlIQg0GU0DxvVpslS3LqxYv6WVOpsPxAX6YpfgsKtUKiup
m8UgnZBgj6FkdiyZ4l17pF3M3t4qVikXvZw9RdDUYqjX2HYbe6mHhD91LfXqgKN4Df3e+vWWB1CW
VffX9dEkatRoG/2vYb5VmrVBnVTaaBHBY/g7Spvkm94UqxKzg+KCjFbfuuGPKPXxaVbiecRWWDoP
J2SfN14tdSb7nM8NYfOJ3/LuJ7iejmkmDEL82jzDmyATNYdsP5y4VG8CL5FhdTmjeuV72Po/MUlm
nTitJIzZ0i2orZKQ7gLtq3lyZnSZYZjvp6xT2docjObfQkIlkW6rdUDljhPYM9jxF08q+PSqOap9
SEvIzTyYFP3hqD0/oV+Sudzi4VWpvB17L/BGZY/8mrozawvaZuyEblb/Ma/hliahtUM3/Du4med3
cjo6dwwcHPdrc117wdV+BiGSn8Dt3CGtrhLcFkCBmQtFGMD0Iq4oCd4QKlCl0JxA5Hmqca2ffVZ4
l38aKy2jKMPKkywXg+WdrrL/vTVEJO9C1y3/gx8nqKuW97ELNQIKjaUVBc2d4p8OSxp8wT9w5/DA
XfHK4pRcsx05FTbk3vwBkp+LfNkk0xM33ZrvB0YfEqQLeSRGuSEv8OHJbmq/rm8X0fyw7caAB3fA
H1iBknXlTm8oQm0pBwT2zqjRSDAdXL9VpcGi7tn+yDtNt8QH1YoyhUASN7zxDH54O195pArlEpb2
9Zfcy4BVwt3n1nkDuXjHmO5hf8/jB2nHLYpxiUqkCOyay7SKdCE2oX64idRs19Yl82LW0jjbZXSf
Tg5vNe8etEp/LC8FRN53mVaSEJJ+bab9t+G2PQHcqMQAtzOwjzEBcfCkbif0cdJbNYwFmtY++inW
MRNWLuf8gcwAUqBkB/Q9WViLBQhBE7bOS1EGGelh8T5OFXki2PT4DfUhGRzd+0gvWGO45mvgnunB
f6VFiU6/lH+IwXUEvZOiFy8Qlge1RCUK5LkRhxhqw/LxGAeB/RSFD8BYpAYTxM3jQIFynbDV+HnM
bgfMJoLF4S9j8y6mmPYEqIp1J5jg9PGt7dlYR7IDFSQphg2MHHsPSLDcuFwI3dQKvTcRmlEqBew4
mBcMIWzLm5bCELFiDixY7P1uU0PsjcNxPAPAdidequ8tfHaSrZZ4oJT7Nn2xEJchHrsw2bKfy7mq
l0vOCBAhG1YFv+dppNCO0ErBkfZhIR1R/zYK6EZwhD/rI6b8ZikFjcySvfxMHFydlI3yZ7E/YN1L
8z1RKyPkQgJGcBKyodgBmvv85hrm3AHDdMmg9XvXyZ59eSb2t8Nr1xHvYklCN6tc3oBve3MyWxOj
5ivH5zT3YEqVYesJoi4BDrP3IN3hweUYYNFWkyloKkATaTZcIf/4Tvb5mV5IgabvmHpDt5rPFEoq
U/lJJVtehitTMMtt473e+TieDaQ8mSzBMsfgaXCfZJcsXzz24HQ6TFSWjzLhSKla3U4JsLcr7MmV
hsOD4rqkujvs2M9H3AEAV3TITWMwNWFbaUwaZZ/cBSxIWEuC9DY7jKlbiiMviw1i5suGuu3Pc1m+
nJE5MiqCO6jP/PsYXc264b+FUoTt5wrJ65pka+32klanneSvotbD3EZBiajCJ5gddYJuzRqDFL9M
nhVvggwBg1GhpQ2Cac+By18/WDn1De0N3x0pFCXJmG+Hn3Kno90x/k5e+JzNCTDqlvNa10TWcb8K
s8nHum9PI0EARO+ByiAK1wDfv0HuqLbzJtnYU2roBcsLik1i8S8yjTUfae/1wlOZSOx359r5dFFA
t0PqYbbPBU0wrDnng8T16de8f0yMUyZlEOuFK7twlv0ZxNQiDaHXE67+rt2OKiF1E79q8rM8n2LK
Ou0AnoNwdbS4LVC6ei1a/56+Sx7BTL5PVSZsRk2AfpQ4zi0CKTQC9m4y3eSXDJNWX6jq+wQU/MDP
gUfPRWs4twBER7giaHQCl4IooTMdsqdM2ulDsyiMl7nLEYJ/1Yve/+abzieIKUW3dss9DVwTHhxV
/hNv3e440K7o7oxX9xClKhVggoy6ydya3U1bwZxv7feYsBmdEo44chTS5plBOSaNG/MluphHh3s8
f3gZbJUjwBXIYwXQ8x8J2KQF/C5oAGEjtGr+gXfRmmLq20DeGswqkaoFY0sxWH5acepHkFWWLm1z
N4+wBei1sePqyts5OgNMekvJ+AyIi7RmOGrN7nlXaIEE26q9c8TYcncIfnrc73G/FnMAiqN5e04h
6KcVY4wt37DaaGMix7l4alL2uepnOWdR2tPf8FgdvmCHLeOZp/5+u/zWe2OmqfmYRqmyKN+kOy/p
/gxdc3UCjyeKi4mFlhQaQiAO9wjIULILwbd8i/LBY5OBKzx4ytUEMc2EMydrZY0WIUwrVqxBllEN
EJWo5AFkfEd9dA5LONYT2CANr1RGl7Vw9GR4chYPkxESItTWl4ceLLp4pD06+J9s46VdUj/ObTdw
Ei36uNfTwKIrDy69Jnpzju39h69gh1A9IZ2/HeWBAO0thsgu55Vuzuh5mnc0Sc0lzM5eyPgcgjsI
IZrF3qBHFdA0EiDEzpI1Py/9Y3vlZZNOLDDAulT2gjFMxTIDsROBtEvADK9gyeX+KDAmDHtd72Yz
W8gXdIXm7goriY/vmgCmg+C2LQQ9k8Dw31a76873Ftw+G3/RqF2cnSXSCoE0NYO/qpMQN+j5ecf3
Qdt40j+6MMYmVhpaQGOm6FPOHCPlOrlPQ7LsfIPT++e0iRSGG8RHY2AgHR4HDPH7zUj4o2c0lMU8
J4XX4cZnXNV+nDuya/7pTnB1ZTqI9669rrQO7PDgRd/lTn873wLYheGzqzW9qY7A8oAZ7jbYuS+o
U6u+cb1H78tP4ZNs3yrihvMA8Qn3+8aV10MatSnt+Xsnb9sDXoqTmaB/TN0B7AFyM1lYwoZFQL0D
muK6c6xjzRutxKo8YxLGm+za3sx1iarU75WJHoAsZ2LmA4fSIZvpTwXrjE7IZ0P+B91pQcAvRH5s
LzL0kXznCwxKMhmSkzDydpUACsg8B3Op3LfbaOFjY7BvqnhT6urYDlNFM5n9rsEkUKPHJWHSpwD5
v3ik+PJwEioR/1McjzTxo0x0cuZNO3NDcoZwLw9agKAXG2DG4A2SPkAD/5F1OB1jQhvYQc0h4s+d
62WcPJ/1voAVGimmWJMZ+9VIrUygRKoaR4SwJrYMcIvChAz1AnxiPK3giuDgqDMZYnNvWV1oho+r
BSqIc+OSqD3sVHxh8AARjjYaLmAihUPAgYDdLcKY50cPGD6MnPHdqoH6kTBhojAAwbv9+Ax2lBN2
j6cN7+ViZT+WgMLlsqPQmYulNb5YVcOXZ+0+0yoVUNxTTeC9i1qdiKK86Gf/4bLXnPk/DveJFLlf
S3WcuUMtJ/mDE1Z1+Sv9E1WViCtBcShF++3Zv2fl+kNZDu4GIw0xsynwVGQB43xETq6fnp+oSSj/
Zol8Lvq5DGVDZeGMZQ45NkzI5SMqcasNCZRZdeHIWG16lqPFPVcibT6x8RqsljuuMTdH6mKVzoVw
z4mnRtqTjC0YQqPcGUX0HS0jGHhGAdCrHqHu0k3xCwhw55tP26cquWsn9fzxOYAGPLfTeD2sPZMe
EppDIoLpoWD8pa+BF6jw7gLvrc2IIiZfJjHYGimcRbb9aRl651Rj/Q/jwLnK/2KzfE5x6yDGL7XS
tuEkux/F2E3Tm2oC4rCgbMNSl9VKnaxvysGmEpaH6vwvUaVgL4Rlj9b/9pJ8XzVILRWoJoUeVUKh
wSe0p4uKJ0Xw9ZCAgY/tUZZ5BEkMTvBICJkNGtZlqhbTZ4ghUlnStqDRkayhgnFciZEyBXv3u2c1
Xh3zH0WrFe9TUjHIr6RCQQW6tkVrq03CQ3ZC7ccu6TJJpWPNU8uLyixLTxr2EKwNTPWWpy2dB9qo
yO4aaPMMDiqeWHpw0SKMZqUCHITKVQeAYDCqexVMdtxTTGXnVV0dKOcKFVaqq3Fa4ttywDoQBg/R
hiPl9sDBXaTTNXKefHp2PoSuE/Qnj251pCO++O+h3p9r4Pm6J4+lZDAosU26aWbvMjHBv33Z4cQo
TO8I3iV+9axSWaLAfAWImWplF6Tw+0cOR+5zJYYzaARjBZlBM2ytpYRjo1Gnpr7gAFpwIWpx1kW6
WdDShHnR4beeI1EtiybeLQlA/iOnypvZszQrO2K8xwUNrlbatrkmARtI5A6Rop/wuf3DE33PtNZI
XRPpS93tGLCRTa69lhZF0YUppYguc9OKg3qeIUUiRaCTNEI24IMwjVUftf7h2ubjuZ0bLLqpXNIY
67kFdyRwwGuzxjjEA9E6zxMKe9ey9fL37Y44pbMYSQ+B/PCtiwQfBNmKgdoDLwEvdPoVKjQh8Y2R
24AIDQRszvAsToCCkXDX/AmJUbCoiq1xe9zmA9cI+isY/l71TPhmadKegAknoirOfx/KRfQB1Y79
NtyyxMgUu1A76c2wK04JDROZUvIYhqJTVktk6WqKEiDdhS3S5XYxEqkk1/nIAU44K0mkRuFDTmrg
FOq9ySHRCMd4QxUFSUgj7QOW+2fU4ST1Na52zzeBbTVKAH/YlffBfNKPFNV9nByNFxteh3ZBUkLl
nfmWNrAh9XDnsXd5yjzHN4/sL+QILjK7zklxUfoejH+Xlrz+bFM5/ZdS8KhoJjcBk7Da+EzMO3gb
7aR1pkt5rkTZkMXaKgHAKLBGmIkJbOyyPGa3XGYmWirOXScSjz8Y9uNf2SehPimDTzLsJOckeaNH
SOLjzQzUtAHi7GrtN9z22oJVPk/OE8eciizskHW6IigTsZYqbuQI4ZlwxPUJX9ycOF4tAaqqDxsJ
+yKn4AxbgH5QnIA3+og9fMGoSQb9p9UX0BpWrgtytBmRP61+vxFjNsENFtjSPbF6sWZ4XkEjmTVT
Y7gZ4K3gwg73zdWH8BjVbdYbG8gVWI5MbQJ62t0CHwn7nKRb1zaOXG1hyTvDf1HxM2ky0eTJNt+U
vU1BQ+0qRF2dsv0qGNACnyLSZO4OZRzPadlWalIq79Iv7BZdxXBLk/u1KcSm+U4hWybXxHjSwxaT
vvBV1/8saI/CkLFvdtnAtOoaWn1x9HuThzixj7K44JGRdaAQ0JzPMuKOBILYKRDWVOSKiL/pkGWM
lwPDrnu624JPgSkBA6q4557irViwEdW0WDnl2Z11JLIZSI+NDdF3Z/JV87lMYdnokTJnPQdigvfD
CxQOt+Lo/VKAW4GBvCIjImssG8TgTA2UlkbgFD4MRascPUot2vRfsPQhPivYhpFAYZd0t1Y7B9BA
a6F/3HLG/BBR5i787wRo17upGLkRRpMQ89s/zZW3lmuivORBVNWkhFRY5gTzp8kAN/KCVePO0eY7
QQxksXpu0DSWJjMrwp5BKwOjkPkXwELqW4esWV41RkQatqmjKuFd867utLZ3gVh7goEoZK9AnY91
nOhy+9Nsb35gjAl6/pXzKrTlJ5iD77gKXazaM8o62DqhgboQsovADJCqOIMd7Lu2okwlyJTzVa56
U+UyeEHtOzrgRbMXpgb1gUMuX36x8nxyILWNEF98yECFSx9KpqCD91ixroqLMmP7HKh2n4TO3hI/
S7/w+ELQClQ9bsAoB/6UxHQjs54MNrERlo/l1HxD+kXXxaQYbDUcvToknUneKejQbhKmdzB+LeEX
O+cHwsOvI8xoNalrVxGS+pAAlVv8duwEg5BTXUA2tsmPkPhU+j8FDyeKzVWh9F7R7qoH28tOQwIF
f04VGLNEpaRXSb1EbgczSuGvUZsHV65kdNtP4PoswyrXbKQOoCcjqcqmi2GdLXzJZ0iQWvQzxBBW
Q5MI/cFEdcdAzQK+j8yc3YDz7VYMiD+1fOpu+9ryAIkBrwJ7gPHaHtj0LVbhZbHTiSFzeyoDMGoR
2nk3w0e2uNyBl5hJSYwzkgtw0FdmacvSkxeR7GA3+phkrqVf+9Nmwra6z8AdhHBOHmTFViTxzl2y
LPcqeEocLrF3M1nvX8Jwp0l2EVZ8WJPSQb6RGT3J82pWFvnffAXByc75oox8rDGcGA5/a0Xb/ZE7
SF/aZYbjA9yDb+IoMgn2LQBsMFHij4duWpdPJ77bS6H9DZNNQjGD/9QzLODDvfvzlpd3E3vr7UeI
0OKyNijiZli9lIAjdonhNkRPsNtphUi9qV3I1BjvzdOyG4me6R4398/qoR0Ua8+ya4GD23G1/iXn
zrh4kdXPQLht1DUgJHSADTn9cfnDUcVG30rX6LAxeluPXsrKAASC3JNLRowHpQmOK/I6K7BySdlX
m0oYifWcddrwWHBHf9RXS/8L0g4AoYd6wLvhruMTRiExJBAzbcRHlBOYu4ZvfiuLie0copvcf3gc
qzLSZi8KpzjgbUdWonmKPjo3cqMHDVJX16Kxa/zcg76VzF14I3728cf0nvLsdYKT4bxZXZWoLfXJ
LAtdrdGAudaOYDPE052OwPRqcdMLZapQRdJPIvdqZsGr50WikDgXmZeCWqs2KRR2asLegIWdx9rz
2q2839ibSSQfY8e5v4erl16WDRCM5mZAgJy7Q9bt6NNR0qXjVABy1J2ksruEm/am+l+okMYOTLDy
353jbBRyJ5Id266JYfghQfutiz0Kr918H/Z/DWx31c/Mhwj/0GyOgFpiNcVZOTN7l6hR2n3DQ5ox
3tMUeQ9/mOafmOcRGCqyHKdmdT0xC1ybKOtRF/WJmF2FGVgvc1BhgGVXkTHcAwCNqHiujxpO3+Bp
BU1ucQbMGfC6MwLJ1pJVfEN/3irh8eoiGeZgJPMBRm8Lc9z98PXanhBnGbJ1B8FiA7GqT88oODlj
8mxXjdgwXr71gPrexq2CYe0dY2gFvIyIXBUX/Mm1axzVLgLteNiaD6T/2oTfh7a3l9EwaVPlunAo
fVhXr+R2M7Hsg6cWH5MqfbJO3jizOBRlrCcSZ+T7Ne1abqMRk0M+6rDLpv4W5DpjppI1WpIgKjsh
6zKISmc36ibL2OKmZ9rDfKt2I/TYO0kRy9e8AW8q6ah15bICe1kU7SSZ63BRLiQySBTwQwijy5S/
cszKkII/ETH6ZFxpPKw177zXAHDrGK2IUJgzN9ZegP2S372bDDrDFx9TFVPjE/iweVO9a3dVai4l
uafPpuCORGh8d0aZkbznRFXsXWUEkia+212lzOBlf1jkZSHhwnMIYs77oH2VyV9ZpDp61Nusn35C
M9ETNtIMdtbsdisHXwZo4wl2/Dwx3EzjFR8YN0zDSfuNnBSdglTsfYbwzQEgPjfr8GxIUDb/zWov
xSadKb/n4YE/bCxCmHwFzmewD1fmzH+ze/OprcjNDnULtgJ2wZNx1oy8GDUiOeeStE5RUZke96jk
CADkR14mTqUMC7ngfmeP+Ekj7CjKw8s1XEdOkktbMxMFsICuQycevnH4TJjrkOqmTPBL4US5nF0d
Iw9dWCR0chrhymJS9/u6Yd/KDx1GzFkGR1Yl9M/p73enjbzpODJXlI8kb78TrVIJe3g90xFf/Z6i
zb23SGW0PrBw+7Rndsu9Fxp5sS3g8hSVdW2b0fYH8bZcghJ+CTGUU6alrivOX56MV9g96T+OguSd
e/KqT3ymPz7QNYT5/WqTyCLmvtNFp6u6d2BT0SDnflXaVk2o1G/MBh+4WUsXdoXkuunb5FscHhb3
2pqcQtNBHXHStz7GjBTeJF6ONfKCQbTO5Xn9MRdJrJv1umVQ5iA4mJxGVQCEGoH4AHqyLCcNQWAI
EhPBFK6QrIDPLyL7N98gqrmZB55Vv7GAwxb1ZoM5pArhaDUI3K9jTTsv1ITye2vljieizc49NqZY
S+W2wSRXow/4XojT2xKeCIkd/ED8gMV6rmWiDusV+ENUB5yWHU+q+07ONJizWnsNdlxgOiwsMkEC
1pqgd/S98DE7PBdAdg+ov7+o5vZ3fHKTx6h15XwNptjAKG69Gl+MJzFzSlFOtHqUohUtCfXr8rFt
v9fTE5ajv9Q/OqsWqNbnFIbnOw5UqXB9T/yWMrZ4qQqCiqoNigI7rA/NFd6VWlbm1wGcRu8tCBJW
SE6czctfNXwDBavLSZ9ma5k8eyJrSAiv62VQBPns7OOHo8OVLTiJQ/YBmuxtB1dR2sHiPxyfNbZE
RZrkpO8QlOB3KDIcvmAeG2YhPKvp8fCVeWgjzoV5wspnwJirvO2gav14KvdDbCf8iAOGYiOoMdMf
beftKsK3yeLaitOIgqKkxaNhmnD6OOlzaFvZzg0inLDpr8WvfMqSmaOrytkvE0/9wGmZiymU9pM7
dO570eDVJI+kuYOTo2vhW1IGFFt8h8VEe6ZlPmSEH+M6OAJTkHOUMBNn4QVuPhdFTMGGajt69fCM
IfhDypzKFtyMCxZx4Wih9PL0uj4r9PSkQq/Sb2FkcS3zBkRaQberpvSF8Z+TeC/JCwerSsBSq0t2
wKopaYpaLIaKQnMpQ33Nlo+Y2w7SpA9NLMPe0uU0UDAU2cPqBgup+AozEcOzG7CCh0BlC1Mc7EeM
I57MTRT1tW36b2Zf1MMhpdSQ2YgFiFJjsdLvzMW90EnidK8jI3RAaH5PQunNVj6IKIbssgBpsV7Z
GGuOVDvx+zxJXtiTfx1NCAprLuo31X+iHdJdTiXX/k9xZLFTBuiugvOWrK9r+la0Vi8Ygc7gEmiE
h9U0f4gkxlqhQTyZiMg+vmg5sxel8QvufGdQsxjbKBY9Yjh9Lt8Rd7KBETaDyJOeGligv82Qyf4x
Kk7SvLp4ycZl1JwbGC+T+fZf52EUte3Fi2qeC6CZS9abrJ4kKQBlZsEi+1RtL+iTPs8G4MLQPeNy
+7m9ggRBFGI//MIf7CziA8qt9Gz3JeDeI+Fgf/SK+fvRBv5CY9DZMG8x4x1Gwk63lpWCPXT/zT2S
PX+VimvFP+tgSvTd+2G91Ah/4uLaRS+UDtUsPfbnIPgk+PzdJEWS8ypUSi/yh058rocjatSusDRT
939ueYwOXPbltXSAMWFUS5mGKSJrOD3N1F1B45xciA21tSkjdMdhBhXcA3EuZ7fKRwcC6mRXyIvn
LNfnTUMkbSQn8nqJ059VT094/R9TDKQbFShlbIhVQ5TsWDYquSSaOaxbS1byf/Tsejw8S0/4S/tg
i/PK97l4/jMvy4WG33yjB75PQSjAkTvB7hVL7Ksdt9B007LBM6muHTghbOP3mXFS/XOURzuaNLEx
+iKBY3GqtkmBq4B9s7VDJSYAbogW6aW1EaevLEb3jmxHO+VDrrsnWTExPqu2TF+D2cpkSmyua1g1
Cl4WQzb9lqur9lcTGysHU7PmVT1pU02hHZEYDlIDmpSJGar/YUg36vIgFHOrn1hfUA/lEkftUyqt
wgjraAUMKvqQun99WJ7FIUnshJ1PrsWKu2slA1VHeTTwNTNL0ylEn9bhcgAseBYqR4YN8lAFkmvz
VLh4KFKM0vTUVol6LJtwpvwtUCaQg51r8Fhfy5penxuoVOpGIKI4S2KAFd+kBBxxrpDxLtXlEONt
XCb/oQlH5SK6zzTg62ZXnEdkfq9UAjY+D79iQZpl/bSbJmBeuxZUMvvs/N9aLnRdTy+/s+JAKVoA
2J/LSoMFCGaGrXZy1XBzCEa8HChUXNImppVZ/VLCGaDdeQAG1pJg4KoR9ChEKZ8mS8p2t0XNVBRm
zvkUacVpXWfyeh4QAs7jjCROVZxZUaIgy1iFwkZLYLTxI1FcHbW5y7ZISrP5Fv3s+aQLKbi2A2c0
YOHZApGuhAuyCxyCbVxmFtWw24k+0D1NdbclWVAWwMLq6kGjKrMVBE5kintYMkd+ZTdq/pRO3eTV
OwbBhl87QDJmcgchMYU1HRvRtyv03gFjdjWlMPg5wlEkU3SDjAgyUZXhxz6r1vr5KrCRQIdYKKRg
8TVzS3+VK9vuSmWaXTvIMKMPdfTRVZkqkQwzaSGlPXKn9GBmJ8DRGqstLNkUkZCg/FOHqoKmPaNM
4AD2HaVb8+4kNEb4Zy+U2+GuF4UghXxNbe+lpPrhtZLkfe+WZcWI191JjpYqG+B1R+/hbBm5p7jd
avWVKtfaR4I3FM4eNTcVkRVsLzVt5VZ/Z4qs7Qf7UuDe3e7jyz5mS6xVlobkI9EYcpeCTab3it/3
IGNMbxom2Ac8hLwy+ieKYtInK64PHBMnrasoFuJAE/7TJdBBMF0je3xvHqlIJW6VVK4XWHmIWyf3
PoNRQfAabzP2UXSfGoEd2d8tPpwMbZ1CybhFYtK5XQVObvgj1U3MGPOGHLh+I6pYvsLuAdk6wgUo
TyjCOEdy2DoTiuHctwKT3GL2c/vcULQ/w9eobk/q9GzNkLEkMLPJ5Wy0595OOjiakp56P7bA0GZT
X3b/VfsjVCxDlMMdopCbKo7efqC1Vape15CHd0rBVztWuPxg3fwup7bpaJdj3BeCFWYTlWLihbk2
adtK25TI9K/npBe6hIw3/w5Rea1IrXMma64J2OwshJPvnIZbLXkuVDeJadSdDzAydEEQpend6rXA
ffOH0U1YuSWkNbSMzivrTUFkcAKtsPiA9isoIRRTY0xhOjPz+iueKB7QR6/429NWCdpnNKjoWzkH
7eHR/CtgrQZGZRE24Zzv7ZWvI8Dcd1xX03R5wj3XOd0QOSRKYOCb+slKMJ0lEQslLgche5r2qvFn
wW8CXpV+MjBTUFtC33bMCCTE6JEx6+B1DtNScV3cjKcLvoseCis0Q52hfugbuTMKva94Qsj+0uUU
KeOvFgKdRu/ipwOMS7r8FiYC0y37sXN7MMvYoanGIvsHPxBqGsx1JvCNe+p3DHE/s4uJrWsHlIDh
Je+BRMOj95LR+q18rx7fwe3R1f5aIt5q2vqBHKb+KTO6chn2fR6uod8Ufgi9LP05fTqbfV3eoD/7
wxDWPegS45sraeR5Zv30q2v0E02EKucWxP1nWsnlQKrZdJu69bgzbEV4xCWEuycNuzDFFIIZ1Axv
uAOTDQerHO2AN7m/wNpoc7LUd4pjMj07stlAeuq5FfCqFeWxZetHnS83BkG83VgJKS+IwWycmywp
NwKsGAMAdDY5AmpUIWZ2ZQtgTb/F5EEIWDcD3VuDig0Uiq2BFnXFQARi/lNHpyGSFKp6NNA98IaR
N3A9dFxn2yoSwEOI48ceBY0EcDd7vvGFKUfA3AVif6lTrRixuQjvU06qatAQbZkVWXsKXQhIBwnZ
pvB3511bKQaGk+S1djGTZ2+32ZB5zHcdYJscP8r02pF37nyaUQaRqDgNRbGSs83aeW2JcT/ejMXA
TdYiNTHMnhh/yETH8JvfE22DEGRxyzSh7niVERwHr9mkC5OeHEqHkLCwwv4t8LnPli/eKHyWYojy
mpmwNVVRZS1jQTKmZ8e/7l3lSgxnHZHaDhInaW583zHxYEwBaaQxhMSseGlUES4lwJ8cd6N+ZykI
+xwXW63929vzejTgv9WNKPV37VmdrEoNQWgbuXG48JYOebxNOM24Et/iEODbfbKarBcpUVLnUydY
3k5e4vTUMQuUcEpqORXmhl2D1COtB3WMgGC1p42FwshiLOseLa0ex/bgsaEb6ljHkqQpJWtTshdA
m+BrUPckOD61Ccw7/uADmdx2eiccdWahCc1k3s6/0vQzT7zgQmTGo0IfoIjv0O+rv4/lwwOXZHxe
Yv9rgAoaCbeGZHerd7hD//1e8vk6DWddrvi8EgnrQWwaGL+bAW9zmSxKIltY+byJlHr5JiZYXlFO
3nESreUhckOBWUbXaO7tABp656qAD2lNivMUXqYPBGwg3aVcOe79j3nOkT9UpWFLZcloM7cxFh0V
p4zvkVej8atI595vsmfCpqqNrZM4SSb1ksVlftIYyHAGsA+PGFRc+SETGF/QWFmo/je/NYmasLQk
SQvSfyZDN6c2UwXjqieTqWKfDeFAX8UO4sTTGH7K3UUtcdwiet03wQiCLv8kne3Ow71if66u1jMK
QLWtyXMfY/wCYwvZboTFlQ5eVFM134jFcrRQGdEbyqxujFGnnCPalCTggBYuu8anYeiAhanoAWW0
qMOrsKs4HUnySRCehIIlsHi91ONdMdJX4YtOAgwii+lz0Um+GX2GIJS6j4PEznd9KolE6Xk8ZYtF
HWccR/WEIxBSG6Fr4McNbHbPOC0Gjxz/SKzoJV/tlj5g9l+OQ8LQ2xfXlerPfw6ybtjxPKRQzN7O
vno5BNkcsd3/DEPW0TQqbyoZL5Bj+G93QR/nwFvTWIyqJ5qnOc+t+JbNurmL64O63ypsGbUqTytP
+MBwYVVpuV3bWNOSzWnxnIum96H31mGj1pLwUjiPRrnGpQrh/mWTDxp2G4X7eKUFdkmBAQUxotbI
7jsSiXI+ZQYBq4DiCMl5a3/JCdRgz24RaeBqCuNow7IcRIDnd56hkRjf2GsHRm1+Ec1bNX5BFlk0
JVzfvQ54Va63fOJAcIQOAK98GFF6YRfABzRCVDHrFb16bny2gjW9leUhVU+PEpy5E4IItL3jhb6I
iNTZE6whTvNgYJ6M2UhYBnM53KLgZJvklsDALhbkNn90qDewKVdwnOEvYgRRaVAOQ7TxfkHu9UPf
oZ8Y0K4gaqMK11eVLY8T+/Yiamw+XhsOtTiOHL1YDn+tS+MjKgh4MuTguJcrCCP8PTBIFrOdkdpV
MiCQ2gjFC/MYfTkQwyZEz7IctpPAVUHExi9yxxhXjUy6wy116dFsBplikuPlt1jy1WQNTn0iygc6
fu4LPGdvjSbZ71TkgQ5VRcIRpFHNgCGuwpoc5sivk353S/s4FnS21f4RKyl1i12rB6KCQhSoEutB
G8YqlHNJH1ySgSi1whd4+zFK3PIEGgDY+jk990xiKcDX4rAsXPz+YBGVyLNkSMr6ySQe+J6xqP8n
BatqCRHOzuqpBfKiacMP0G0yeNc81LG5gmO2TM5kK7mnmQSOjPeqojOMsd5F2mrJUZ3hBrZhIf20
rcMDMNqstTSTEjXOJCiXS/ugm19BdL3VwxUGb4Vl+JKy1lD59THpeZ+g+tuKTIUsYAwvp8hLaXmo
f8K4qytwdA5CgEM+FbLtYJoQs3qbgJR3BVBS6c4bkbW9kTB+HHvcZ882MVh31ZszdGvqJzTczYKI
nQ6HZbsCRsHINDYI4TQPsnoRMBHDyOB4p/Ewrp0rY2C3ZPfAptfLC/eHkDnWAP1OXcW4pkGNSGsB
JY17f0Gm7xJUfc0lbDdtO/ZIqJxsmsEisUXUrtEPiecXCgyAyiNCTq6jZHCaXmgYDTjpn6KD2ZMq
QvZoRfVoq5z2uL9SRojjX463pXCBFdPjL1zWP/SeU7i/nf1nULomN6c3FEh5vyjLu0USx7+cmvaO
6BVeIKf4tVVJVt23hAYss5MaSVepwHdNV4hj5aUYMWVT2vvrB+fK5jSpwfoBF+YFflIU1rQjSsJ9
CDIr33XAg5DOsLRxXoolb2EXzbNugjQRDvUxkB56NvBJLGDGhZW712PBTzq3N4s8NByW0Ec/CO6p
dFOp/DfilemL2LqgnFhxodyboxSNIg4gVCMcJSBqfa00f6tFh0Wsyil+3AovKu1gdiMfAzduchqp
8c275h15w3edsD9WQoecLS7vsXnci5KKXuTzwwBcliy3lRSdr+kfg35lrn1KkCmGgmvPG6ONUypd
ranXlmWENkScrnLiYxg1rtn0+694uPKdJIte/ANwnSE/My6SszC8/eKn7IbfxVLc+FLavz4iHh9C
mKYGuFg+1nfy/821UJ9XKUodcwseV8b1+VyGI2ntSnfKCq+0+mp9HnpWpTX7oaaeSDt0WvNalRCN
3xb+CzmYwaW7617FFpbdmY5s2s7nEL59hDZbwWjD4LRluhGvaVOss0egv9xThTEFyggEyf8BxFkP
ljvJ6dHn7+xtynsV8cXolw5fPrk4SYf1lGUg2m13OWtS09NckKuKhKpMweF/FlgwDsPr6DdiP53f
782QUm2xukTvDH+kwfnMu98TlM0i6D1a0WRPqmSf4HsoOsGWn38oeVfRVuY8zEkCeyuR4H832xU1
PFSSidEuFJdfXT8zN+biLRLEqTi0VFLpyLIuvOG2uuRZGm0gx2ZfTi8y/HUxPp+gCGp0pFbxKULM
8wt5RtOoNBOVCCxbUAQHQQZRSVxBfjqO3ZcCS2tf7OdOC6Wfh71Zo9UGLKvVE1Fb5jImKqgkxLKd
2540t9gws1Qx7KUBMXew6PjIjDLVMdi9O1BC4Jm5PYSH0iMiCz9noRIPuJBR27JxXokdo7uRrmqj
l3B6B26Lc3imTgEHx3KH+kg7ph4Nv2mEMJQ4g94o7BYqevBnikjkKURPwhDVatUdUV8fH2e3W3pZ
CeM6PiKVMYRhkCQrYp5ufOvessTAD4EY73GHTurG/uKYRXrR+stVX5QSiucmNXhdPXu/sQqEc8JB
NUjik2SKRryZXYwvGmZ+Vs7bTvgo4wQStUNxYkppAX82T2MGDkSUNkYZ8oC97qm+JAUbIY0SbqdN
jv1b/UJupdAGvmCfL3S2lkBJqLu1rY8aokawKN7oUq0cuWBkvFqBpJEp2CH7mRAvBUzuRcPrsZhX
gaH/wM871ZPpbHh9b56c7XoAIfzgDbdR5gxT4CshtEPbeZE9M0vI8hs4iPm9kfqCJ2QohRBwAuDe
t9sDfYUubWm1QrN0VlLjO2b/mKOE1uCct0gZ60gG9V04T/gw5TcQOHLJtQHi7rWJ6/JMm143NJ+t
HtSSTGQedIB0cw5/3gxavdGbE/4pYHAyQyTDN+nUj4Eknl+9KXuLQGcrrMYOsSaq+b8N81S+M/Gi
T2tHGMHDoqOk+63A1TANKE4637W3qau38IykEsqGpUkYGpYl9sNyEnnI1AI501QrPRNC1y9YiYg5
6mIjpCtbwxBVilsHdG5HVqQZPd5N7FrJQzQXo39+69JUlE2LMp+YD8DPyV9V4ZM6OsZ0rLyrSrfu
Sd0sofk3V9yfwJ1jdJ9OjnLWS20ScNLvPzg7aIXNc3uipb7JWV6txeIbyQnWEMJs9acTZ+1gA5S1
ZCc7q8YkN8zoMP7uj3KPxQ1L7DwUWgwEp2CMFNd7oXkdtBQFsWQa8e8Gr8EEpfbYNOtrOPe+2c6r
Ss8Ep+9vZL2yuXB+AYN7ZzmTEX/YPn4Fv2NBjSA3Jz6jBo2kUQGJqiUd5sezLxErQ6glggxzfrZ/
7yaO1ER/etRXBHTx0IJxSHwhk8+TLjdOWHZE0pJ696KsZdWfULsQms32I61I7tHT5BGXeXbDGzI9
2QKagfvNzTYs6H5ylKHJRnnUU3q+gvxmCO9e4jMDvVVMEMzBv750n2qLIULCYvUeGOPv+lMgWmIZ
YyWPy/+nsLnmZ7vNOc0ocmzgiTHhlFwNfMWNP53jLH6AZS4rDFpsD6UCEN6hbSq5fCZqioX2FIxG
722WbDBXwW6JJChEMTxViQlSuPVH6a2JVWQ5fmWFWG89FAjpZR5AwIIBn4TavIU/HAnNROg4uE9Q
dw9TnpJmynb7AyQQqWtnYwA78PMrLwqlTWeq0nn9n05m/2W046yqAyaLp9GiJFK1Ufe4XAdgMOBD
yGeImcxAtQc3BrK44O13TArugvZWH5k1IUYqnRbcuofK/+U9aRgUL86DdwTcxptlC1vlkT2foObM
oHVq8HpPdMqU3AEp+1AnqviaZv7QgAvSFYJN4NHytzNLrpUS84DNiz1OJ+4/A+bV+m67SFeGbdaX
DLifC+UnHtnWo7PwBDlu5ROIfOJVz1xcF5xlYexh9y3aTQQiDdpSmjo9PukjNTAQVAMw1lO1tbD0
ZTEtDOBe2mmB5Xv6Fpu9dEU4//ncxwFrIIGQWKebDh8Y97RdvEtx6EDPh/TUBlQEjSCcG/v0cnnf
A65X3my0QBCHtdZr1YnjhJo6lR6QBihoHAkbCKztKRGHo+VRje84vZhgSwSR9yDu7B1NEC03Lj3c
iBioRZyAoJDiqeE3JpLm2eOteqK0hkuAme33fDIe2/A01w9+gP2K6Sq34wdfWaZihkmMY3PE7Sl/
TklrOxFQcsRo9x7mNp1nCZKWhYFx1wIIGHXMEibyjebTw9KRgnIU9IpveAkxdXbgHI3CyNG81nT5
JaEt5vtJ0BggmEpUH8be3xfbUOsxFs+dOwI1haY9qz0QIvUY8eIHNEf72yBDPxtB8Ai9q06mB32r
ob0WAnvicXlyEapwagDk43xvZw89Idfrt1tWgMEZ8HlIk5jRuLdMfeFqKbU/g+gCz0/dJIwiVELI
PnWYQE1m5PemGEo63BD/N72A3QnpqpH8C4lnNXLRJmuPUeJCLHoOrDwxv/Mm/R1RY19FUIljCIAg
iVt5TnoL4mqD0uXkHzCSQFkl9AuwQ8wEK/eQGCYchelPJFg+US1hOJ0zBg8LNl5+2tFa3vw3eNcY
IyOzERc5cO35wZ9/YyvCTxA3kbTel379HifGouI5neQ0f2JfrfJQjg0Gwot16K8Sql1s6+sjhthh
MaKYcrsrWQPeebDQeYIPCL1v0YnS9aSztObLz4Men/VBD/VV/b96WHre1yVAQMbuZBMitx3DLXaq
V8BVp7vlp7nJHz3SRtwAhMueB9iiqLalcDHEym0oVapToLl7nfVYKwTsIAgz1tYqsYCZ2O1Zbmpw
Sd0f4Lsvu3NgyVclzzcZoolKCuEx3HZQp5Uk8YnxJ99m4+XbQTGSOi000dMBmxe9DLF2hpH8hfib
mW7Vhg0rzA5KkTUZGDNmUxjpyqM4TNr7DkmH4VzH9VnMsSZ3QfkbkeVudMaH238mVw+3l2j1vyFa
44udQVS047RfTGStDOJRnMmBLBBiAGg7VuXiUn7gXbBXgV7xVL3R/FwJxM4FBV8mMwGRgIyk0KF8
6VdEdux4x4er0rz7uRnPu/xVaoESfEfWJPfmKhG9PNPcmTK1/vtUug0y9O0yoHz7oqFyv4o9LU+Z
JUSi0Neb7Rgt9dFomSTxx/DKjXeKXoEU673eadW8rSh0C5wlT+lFFpXcfKdhpnAgErSS4WxMbn8I
Q0xTCxZ2Nc+x32aH1a70nQ/Oy8B7OJOmA5xH+wg77sh+l5TOoAPdS/jotoivmY0zHJ4sglG5N0Pv
clf6GVJimy+h5ye0E0jcumv6537l4p/T3nzv9x1i+N8GZ+KiAZMZEvv44N1kV9GCpmSJF3FqlTDm
OSZK9fhntpVUWc4n5ducKDJY+TneIFOAcsdQ4jcuD5stSXb/gixOIULoCIgbNNvDONmUfYubnBbi
X9a5niB7cj6D8IGnzAGFETuTUiCTIChk+kVs3Pe2TrZY5vZt9i391NHmx0OaXaGc5m51kCk+DZ86
H8BAqcq6/cY/24TB5SHUOw2mJl4Jq355DumLg4hocoAiqudCOLFfVUGaSNWJmbR1KBXddPnI/BcH
CswajWaEG6v/JBXrUdSt/zKrUTSc1uGsOGPXCwcGCdgRLlE3l698lMZZrDjYd6oQ2KvWSBpJo9hu
/suGfd5NJBWUFlUDIFZD+ZVzZw96jK69m+lPnCkve/JYSqKOPeVExpf4+SP8j7YfbBqlTWX2dlq6
Rh2AS20pj/oPgysDgpmiW+spjk9cuij3Q5O62NkVKyRn6di9Lv5U3mkg0iVdiE4Se4FL/qnXhE/H
1kFZbpGqVZ5dxMpzCX431rjsSxOEW0SHUkn59BnhiVB7sqxHaGFjPZdr/P1RzB1r+5Jk3h2BOXMH
hW+vyq+eKeLyC/c92cMPW49g4iX8PUf3Gxsn33RXQalCZHBOGi4Iuvh3lngQxRuicsuGfK0BIA8H
HaQKNeGF9F5ToxENaC9dIrk3TTe5NE1cMhI5CTI1RfS7HELpOx66/ifgt+C+btAv+ZqoI971WdUM
oYn2sVNGsI7txLXrJRVbBwYahuaQE9rZKgIzQYb+UWdYn4CfPGPZmpO6NcjTRBpevv28otkdJuGE
jvbtELOeGdcGpBwp6sWZrtHXjGd6w+EMNRbvtm9NJLuhXowFxuzhATWNqV2pFqxov1heGIm1SsiT
5qWcd8Z/xljWGAMq6FVng6EVmg3OjW3cImW3cqYUb34BOXbQCOlHFbbVCza+PGFGdUjVsSlpPGQo
SBIJHuJANxw5xECotoqqkbLgVrWaUYDbA0+jD5BSCE5cTpyQS2UtcEF00vHeDwpqjRxEeAppRic/
cu40RS7x8EO58UxKptf0OTLdWQwKG9+yRYCuwuFqL1DtYJ/Fe+4bRn+Ux7aH/lxLDR9Twz1yW9JR
bV5syDSrKmviJL7LEbSepdGDbexWKcRu5bh5qUCObpK/N4uCZMABGmNSezxD/bypRhEOQpK/rTLS
IzMf2I+cwSvyRTX4ApCa2jYV710QcafhCxPnl+YQFW6zeGGTf86wFMSUrrp2n3xemVIOCf9BR6oQ
kt+Z2uMqpSzGC8BlufYIArjBRlyDW1Tlp+Zz6nvZrjf3+4dYeIY2JDe/xzWCuNNdrWfIhXsuGGjN
Waz+WB7TP+ty68Rq8KAgyTiTRfV9kXLrqc9fnUhHKTdSDpiAcMavQmLiql4S5ajWGBGXCKF5fFrn
bBMoHvh6W/K0K4ZrKV2J68geEAXv9aWSS9nc/gFZqVzhBfygau7817RI9YJWAm2jNxYKCJZC7x/g
raOJPEyLg4bS2ifmMdbIzOqOYzDjY8mrsYzUdsdBv/dvv7/RsDGp9KoeWvRF8wLh6ATfwIuA584U
tiSHducv0FGi6CQFjY0NPtgpnsNb32SgJi9ap55wsrAQr+lzxEypN7x18e9/Kob4kD+Sl92Dedv6
5+by+4PFjSJWtlfXipCbDBezEEOaclJQCm+q3QTwaRkHpErDvGdty488GYg6lXNjzpCwWYAtuTPb
OWZfuWoCMb1Ad+WeL8a6OJjo4kGyQ2efl142wzSlNMpuEueAATY253OlT5mIN81bHGSWO1K08slm
07n0RhKO6Nf9D39HEtbbY5RPTEMpBv2pV2vwFJdKxlukOf4d1Gnhok2AI/IU44sRFI5FRaqGiKxc
r1thZjEzl4JcDvbq8BiE+aX0pnKHeJf8zEewhiRMtw/A8R4bWhZ+5jw626mRO7qN9ClNydNARSUi
Z5EKldXtX2QCQ8G4N7EnlJ3Bm6txfU0SOaTmzqJAKqLZirf8TwQQRWQfAWy04zSuc/uuJejm5f8U
NuE/g/YZ7ASGjUIywsIueAE4A1EoUnz5HRuJAXobhLznuRtFkoz8PPF5fydJgGKL7oBUWaKVnI4/
uV1E3SzCoqVst4JqvR+Nn7m/ob8+SXTGV8pXA2NXZTsARMEoOeBZzrHpvE1IWTmhLC6o2NK9u8Cx
CGVbDAI3pZp6jkGjy3Hv0t1nYMwMyOPgzaV16+IZX+qqYMVVBTUhkxaZWeKnaPmr68xWr0mPiQfF
DU/9EvqZY+nOx8HJ2KvaZaUBxb+Uf3OOWK6H7KvnI073GCYwaoYfsTldJW5YImrNYjwfujMdRkdZ
26IGJFfQWMIHFWBSGLslS8+l7HrSMH+FGknW3dIPTu6Sw/W60Dujq43Mu/MeW0E0S7hjWaiYYmmi
+45xsq26gqF/xBxS1QoI6QSa19QI5JKoz5SbrjXz163QBw3Or+0FHUFCqnhhM2pyFJAufw/BFScP
ySBLm6vSyMNkcPxTMFRld6ftZIwD9z+a86jHkA47B0jCnhdTrHnjuEK9BqFVhYPs+UMFvv5Z2xgo
PlbQVBLmRcbI1eI2eJ+Wz6+TJqZ9idIgdrI+DBwx16FxOcOf5Uf5nyh6lrm+21gWEGfhvXYXEWGw
9njJQwjFZyyK5F+D5O1cHDG7ti0SN3POkGwmWAcaIXT2M/dGlr0A/wvCYsQmzXRxyNf5nBR24/Xg
8Tzn9NkoszJbqCKbQ7XrEKFtJqv/a/3M0r3mxF3vDfqao94Xvdu40iyiZdw2rlGqs+9NSgF8F7LM
/zrD5c+3JidXJxmWYoKuf5aWPbad1T1SccvYJbpnito07wUqtDuyeDhMkE9d8iljNlDQ8O8H9Uxz
xUwQsncb8IAadamPDBtpwl/HtfNhV3MXBG63ESHhyLgHpFAO3w0f6J4WXG01lkpjckwB4j8hsEuf
faLbo6rXnHhgUFcloAaZqk/h0GVQzUhuQnLYZyjg+/ltSozx3Nofern1f585YGODK392Ul9JyPEw
CdU5h1MLASBrD49jm+Xac4Okvo0DPsn3MfcbZafNJXZR1zb7KG9+RXLde3jQQF0sJNZjoZbHG9V3
UfTIOMii9ufjGtiMunDKs28AaIK7WEs9JwxyYM07yJBMCQKStF/oFxoMc7Gdji3XEONQOrmjW4Cr
PALNgivY1BgquK24DiCY0ZHGFhvaJXQYCQA2+2JeIZjx/j0MvyxnhH0grQigavrf1Is4y+PMxpil
ASaJuftJZ6wrQDxewd1hob43DzWVzzX9TfMF7M18JfVkC81VKDbUMxamKIB+tFD+PsY5S6tmMml9
wc/gxq+xFjhqIXbZ+m2K3CbPeAHcb8PpHgChAGfO3Fx7HY0QxlUELBWN4HnUmw+SMCs11SjsqfAW
ZKdESZ0gyr7lbd2Tul1pPZpwccFMJE2OEuNTIAjjQcu9X9veS5rshZxM2GywSYKp8VWICkFCHCm7
Bf7xQapZjl8gQVx5rIpVSKwNMZOLA/QuKa4DMD9uXd7BFnmrID1zaRFhdsIafuRJ38V98NJWb39N
woETZnKo5kLEdtVglDHXWRROxfURucsgOO50eNjx5+zhAsVTc4S60m9yebF/z39Yyzj7Ocf9Kb2f
IPkoBJcsfTx0QzrBU1ke1Mu6UpntXwdbP1WOjYHsfeQRPvyZWWxM09c5+CcHDo7hph20Rp6klo5H
7/H+hpyzDci8GyfoQ6DDyJFb3pIG9aUbUEBrGZWLmojMbbPR/+LHWxHJA8/XT+iPXVCdxMljqOa2
wblyM3yV2XQKxqVnqhKtVz5xxUw7GgRZmAdXGO0FEO5HL0hYCImcpC4jZJl4SkYBnBwndY9CtTHO
l8m/RCyoECC+dUTkIZFdVwr/Ez3PgpUfhlqE0jzG9q+LHY1F4EO/iGXr4d47dInOB1Dt6Qvvu7/C
J+3k16kl5GLYDK6Z2FH3lIIOSsSNVZAmdOGFBVko7mTunH5KRT+I9I3iVPUUblCcW7HQE9Wf01Ds
AaRuk3i03H3luNGngmHT/ZeSMvBtyHsCVZb/2n2ICVxZbgYH+drOnrgl3fZZJ/KIPyYKoGqt19t2
q10+CrlxCOn5DwdODdE+2kxFRg/xNjgaszUhCX+q/DltrIw9BuVH6HM2Coy24nsQLd/LrCoipKi6
Tai3XjlbGcs+R2IpYak09ahwgJ6jnFNdhHuqR8xgtfUVWzzm5orov5bY/Ml5vgmrcKTJczwCLzkT
nApcVlb8fYNRipWIPzCuPJxtHdNdqSE73GwSgmCtnU/PzXP68JbLFKO/474fqxKRBosx5Jw5xVPy
mFvoWeyd8DpSuyARCoUmFR5tHOT6fI6AQGb74COiqPVjlPQrB4g4ASW9+WF36bcswsTRsXocbBeL
Cr/SWwMFl5sla660cE7rKmF0d0RVix4tzpe93xjmukuq77QfUE8+PEjws8TioXqDqfIZQliAvZoz
+cSz5t9yg8eXkyAUbSLmU5oxnp5nSSOJyVls3RN6CXzz+yUapUjxlnjfcVPFvFZ2Nw59l0uICWMs
nezHjZW97n1kTkJMadB06YsD86GDk9ZJw1vwA2JRcmNqSWYj0dJyC1WTcPSY7cTLLjgJyk6ITsnB
xAmWEKF1q3Luw754vF60STYYMTar0Ao+v/3e/BUzSxvl1tVqIx1SfK4BAhKndASHoyynA8HQTNWm
fMvajQQeNbK92tY3C+XZKrzLJUIFzCJRQWHbjQQ/Weh2zxu/OOhtctaeUABtXhvVeV/LZh8hXZO8
X3B5WX+IrDGHxaRZ8jRMW1QsIjT3D9WHRJAddLHiPxo0gmqSk9XOKV3w6GYuwRz4iWVLQZBALtx4
qwugVM72FNgTwjb95u5Z9xvmRgMrOGVXxvvACEu9XxZV+kSGXITQYj2Pl0wB6mAlZ02eEkfgIr/y
phwgxE0+UU7RDb8JzgrsUReIExPAARXQQQ+JTFcweucwUpBVXRjmWRKjbEHR1TLwpFFXQpUFQ7GP
OVlBLVsMrXuRyFZdbidHfAo2S+CNawa0heEKhEtoMksXYb92thZVk2BT/TC454rxoUw5RySfP9kN
g/UsJTaol6A18mIuxKW7qcCebJpw5dC+dIrqaL1wMg4s7fzQ4E3mJEujOg1ricIP8qqwFZKYmTuh
ZdLW8ABHhTDov6LkEcXYS5Pf1twMgoiE7uw8QJJ40gsTTfk6/ATtJWoLlfGuAU+NMtjY+xKwk3Ck
apV8qRh3qxHCWWzYP/D7oCMWLwINnhtQd+czvzGq+hcnVuhTjfXp5XtkwKGj/JZFTwm/6LvLE089
66MvKEyRDupSSvGmuURz3XCMt4Hv4kjLbWUJIydnmRkgPClc1py8tALOC+qwT/pgI8No85AsUS/M
VD4Essh8WoIxMAR1HFZf7MgXEQYSmQbrA/soQzp1lYv0K5FqAmm0+pJMZAb6ki/JPc2N8aaRPMrA
sP1bT/yVO9LnoUj8b9diU4yCQdgtSFxK2Il2xYhilyRYvwVI5Cc0Mu8GENA631QQeH7ZEgHT1SLO
DRPYkT7clrTRKkV3HP02IDMr6w/ViWCjmenuasrY1Oywqr9/G2Oxxll0doGH1MfFv7IkdQng2/x8
mxWb9QLPy4pLeDzkZVGUIHXoFSxprJyXxL8hLzXyf/+mPu9GSCiKl3TmEuUfXJLOGkMosUbfO4bT
s9AihdbLvgX/y15S8j6SYzhHdVMpftFmVXm5rZcWBbpjTap6P0M0/Qk0FXz8bIgAGXhnvqvhlOmL
axyHRztmmDNOLfOa+yC9B62Ku+64oeZEOHjHMcVilKOL5ind8CbxF+Sx4fu2jh3OlY7TXvbjPyGC
oj+Knh/aSatZfuobHUHpX5WhcXX7ir/bSv7f7T+7WdlDKVhNbG4EQNGW1dn3cBVF/WHhGcF+onr8
pjdpxGi+PVSeyZOhL41SOWen+ARUDKGAX42gdva5th6OAQ8P/syEU3o1MJm465+2xwUkSJZUFInF
uBfEANobE2ZSrbIIqowvqY4o03a1OWaT0IcC79SLPgC3maGb9bvSzCtw65cpYwwO9UCVVoQuzt6d
IcAOSZAOw4SrO15zoYVZw2c4ymhMDuBitvXvficKxIEBrj335FznGO0kXbIJFGor4zjNwo0cW0QA
8qohLforXJSyKsXcdfrNu1yYo8Pd1TQdObJcvWlVUbgpc+6MEjZIGjR2gg8NkKwJ0S4twWbAbwqe
eEV3gpCOcSm20z/9EXSmJH9c9So5drtnrx+K7V6sKA2W4/C0AnL3d26ZHEGsMITqAExQBcLJ6eIf
FIn4JIbXo/gTHwyxu5OHE0dF1QONrRXstArKtS9LfGWQWswfZqESy+K8MXDzSl+0sAO2BKpBuH84
cNSnUMiu6w3XPEAriWQXpbK8dv50odwSgRAdgdQLzaE1/t0lLwa2cUibYouzEwvBPIArmv5JIE2y
ZYEhvmL1hgPfsyq+Nb5JEmC2QGokj+YVJDGGT+VwBk85NGIZ4PBgz9+ryfbriRe8IJM6x2ndG+3t
2lfF2oRDdfKz62vf5QVbB6e5a7GBIEZ4XxRBKHfHCxa0HdsBfk3omCxw+JVI1DQOifIALcKjtkjr
BiaGuwqsGus8Jn2KrkI1VJNv2m5sg6Fyp+k1ylEmZyRWpJuEzL6c708+aFglhpHsH/WfKI3/G91v
OgdoDFpZotVrJoD/4iB409qeZHGT53Yu2Hr7ZJWUWV+pjArAc5Xro/NtD0O6Sh+HMJDJyT5J/+Pw
6SRxXXMRkxQNc5ldKEQOl+uiJ8Y1j6LZhJJ6KFgIj6gg6ox+abOOBVp4e0scjC0FY+tb7M+GnLEq
I3ni6sDHZvsVSEFwN4n4UxGNKzAnUMbczafwjioILHgt0+ggIBUuUH1145RUciaWQpvN8Y4YYxj3
o/9+ajs6LwvvoF4atVN+ZcuiPTpwqk4Qac9i4GnPD8Jvrn7tmxDM3oWYCwGRP/f4hK5YlAw4bpN8
+ZTK/bdc6hjWCerS5EVopiWA9CYEaPGYh6f9fUDFT9r5NcLzSq2ql2bMt9E56Wri0ePktvO7hxoz
wZc8Cm8UxNYbN5AaZnlwq2vO7mtbXeEG9lpHBYsl+jdO+Xa3O7sXSYuiWHmTJiAw+Tw4+Z1dZznd
C+Hp30L1mIEOrmAjoBtjKZKKLn44mfgGXbZcsPMY2OJ/SJ4WpTmDz2YO5/m/dhW8/ajCqa6hdQCN
WrqKnhjlEpEtsJ0Kgbvc3sCYow4o9DJESNFSA/SuLzEuVFwfRcKO8MF9iroCTD1iyqH2pwy6Y/sp
O1TYiUqQ9OUQeDcoP9jORsXUvFIzZ5H30ZYm4cA8PiuyOuzls2LHyi9F3Tmgd/PAIOtqgWGgbxBr
Vw9wAGvCnL2ZhMRNQcOmn6HdkOrpyFVYJrgSXaN5DcP3XQSBnMh8BoJ3ivdfGwE6gWgIwkmM+MuX
+YrxNVEXqDeAziKEAGVNlfXgFNAiherLx3ELX7Y9YwdGsTwtNc8ohn+sgCqf4nqQNkIoa1FV+QFi
uYlBr17BwR74/qIkwgEJeDciUNWtxWgJU0pczniItSQlfiJo3UimOVuFhSU+7IcqIBrDNccQISTu
92S5pQ2cJNw2aBkNMVkSmeslEo1/4s0LfXEHm/vkEd3i5KMHHtOMkiuF80pLcSaxTrANOHSlO3HV
74Qi7wt1fSA/KYIgWIxBrTWAul24HhCg391y6nhycReRWet0vfROOcRyovsy7Beq9fXjzkS6CJOF
NRxs4PYd6YNw0pGxvLEsPUFhvgzXTXRSwT2rJjDI6kXMpNFRg/pKxnpd47Ee4g/xm53DkklphW5w
zewjWnfzy8IFnG99wwlNbMZV0+4FC9nKXKlxRfOU7EWUFCzboIIRpu/+DhmKHzLur4dEsoYIp/5X
q2KXzSBVwLZfRl1aaUNsSuml7RBjsLn2e1ZcPvDO27TnYaguxWMkhwDCheFGF5VIIguI0ni/H21S
+xtW5xbsqYHwNe4lhsCa5yUAI6trASoPCUVhHOVIPXL57EGBCNjK4Eq1pUrov/2jIRKIf93W7Ft/
8n1gH1R5qIX26SMjsbTlw92U7VYevBNAG79ExHOBTlmUnecZkkYsGtehzAFLEoBwv4AsveQtexpM
ZAu5ZZQmMq7mrrZyjW4CjX6+zOlKeUCgdF8u9qUND0ZYK3OMN6atv4C6QmpI6vS4TDkoWBjNabLB
QYWT8JqWDkhGvQj+XmZVpgMpbsrTJKwd2GyYF8d4rB3haVprGz7FP9VdooCVRVxYY5saN0l3L264
Y+kPn+bM8OmNJS/mSM04Mz2mHNYRiqMZFhHNNbe++oqd0cdEjkt4lTewJz+6lx9sK0gUugn7FKYS
MWzoCELTfXUQqDRPFJFFPx4nfKHDh9AnhJBVu6z6jtVG03M4MOc91uBbaJfHJi+mdh18DPaXL4EH
DYPgY36X9CAnBFpDt5QGQRKmI1QpEuRM445RCZvEr47UH3kR95haXX70le0JS3FM3fQNCTVKflPF
pMfkG/tnPJqa3or11sLtr4/H+g+YZcOjRM4qsSODv20tLFoArctNDjPVpyW/drnSwAwGpo6i0lV9
lLJYGENrileWk45vuivA+79leXicFf/za8tDjR6Fjfjuhipb7cQSqiMlLNSPM+H4mVz9w+LFNNUC
J1CWIXzgPfK9rlBNiskhllUPcogvmfcFzZFooPx0ylmV+B1whj7ZfPxLSrnPJI+OZm08QDbDVf40
VIj3fU8LoviJHh36XOLvrRusuWMc/Vveb2VsKsHSqyV+G7EaBG5HRMXvwJcRR4Pe1b/2XUngf2h0
E8u2aJt1kwXzdDwGKZ+G7EaUaMk7KMrIBR0I/b/8wvj/kSGi/sY+c8aHoWM+TmlQzqrXzJtj0+FQ
44/Nrp6LF4+pLqtcK66mXTRkZacOuTxY2Y028Yw1ITMCfMozudK1q4CqK/LzBKtd57f5pow0BXcM
1Bv8jbVyflc7DSV7oz6LTpNJbP4dgr+f9AajNASd6uWHlOt0d+7dKLB7wRQ+YfZKGH54N/n5ffyT
lJaoyjwqtFoTqcGXCVzNw1G2edEbzQ05/xAEPzbGlc/05BzbPzPS/xBmF7xmLXePlypFvt4exfsw
2SZdXttr/WUtiiJhC047/scvR6th4lb5k2Es29+uBYRtWnL4cJQHtFSnT3rcVmwqPe0yhxpjvILo
Y8LFvLtdREfLxTd5mO/YC8///lH84BvDoYeLeYLttKaUiF+SggPACg4kqz/7y1NwuRn3HKln42U5
KE6fibv52TncCAuW3+i/G0002z9mFiNB9gRDk9snp7tCzc3YtKkUTlRsLLFgruRd42lJFxsvFjA+
QXX3eijVIGvXC7Jb+5Pmb6winWoctv6wtTWmiUViF/Bvzn9IeXSqnwLiJqFSJW667MMPjRdv4qis
w93BfCQ78FpgbRl2zhMAuOthEDqdOPdPs9emg+Opehgw6ZPx4tCvCNyt7QR0m+OTOflnNvEnpxMC
i5OHj5wxdoVpDhqUGkmobHqbNmuLtVFSth+ChhcHaRs5x/iV1QOiQAimcPcrl6Cw/scQp/P/juOY
KitTZ4ycGrtMmcxyPXCLeBCGplWPtFM/mqwjx6TdNs68eCfu2cq3xV1wxiBNna7uIjNss0fm0lbD
WbdO28wQN6s8bR/S96ltho5kPEcPVzPoLkS6oVeVpIWwsk4NFRQM8d/izz5Sunh0sI/sMXG/pKfL
6KjphvsGn4c0rw9CmBTJBVG33qhZzwHSxJjtfXMlTimBwrGldxVPBC4p6tD0d0COr7kJL24OVgSw
LUsmkbGWiC3XhmQvlOdfwEv6Yp5uecDJkAUBG7qsBn2WrxvyP73a5YbcdmGeYTxu9BKT1s9udhaY
CtpfXwkRpoZAYUjbBVUmek7LGqADCad4oXf/BU4PCvBzfVq88naGx46rGb1TxOkjLhPUU4N0Lsff
IPbzWSs8DjOZEIlbOJaLLSIMTPuk04P8YSU8myWAIZHYeGNUx3CTSZcnYGL4bNYEffzgyxeD5L+C
/VC3k06MVwDlCK/G37mCW/uQLa8TF/qyirEviZcuf8L1OhGrQB8RgyTFLoq20XIVZweXmGcP6y9u
gKMbokToTj1+2qt+HbN+8I2XmN28AHsj637/a+3Mk2fdAurj4lEuJh021w3GOyVZOItDdq3Sd9h5
kft6Htl0Ri7fyYefOvZQG//fZ9YDSAszdu/6ANTBcZOZcwnMYjFKULmh0fuB6VmBuDWK3aMOnDpn
kZKCR05MbHcQes/QBsvvPWhayFsltHm2IrcifI1M1xNVKBgwV3crP2mgpO+EknShd/NHxLIyxNod
KwEAuKhpLEScMZhNK5i046zZIIiVTGO2CRd4DlnJYalkDESyNCt1qg0+ZT1PD5mJLo63L6PkocHC
vmmn1ReJx2NBTK8vcdblEghGThu+VGuu92GC1hc7oXYrrGO3DcYkGmZThnDELG6asPLRNIrg+ryP
IwOsQHkcrvlVl3oPvTSSoVYw6njkMwo0LY9vc3lGexlPkaiX1fwo0LCz26jYAXFgPbISksKKXnaO
AdAULoOlmnsBJQK6udXd6WpvN5dkwaZ9SjbworoSBiO+gqmJzhFw0zaXtgmTDCMNyq9qxLMFTLlr
pDhDTdUVV1TvsqI4cOD031fN5njTSKFiGRhMBObmjon7PrygYMOahl6n0WeFZFTSAAgznGa7kPZx
R5TVoMhtvcRwxobAt+qeLMKw56Uiql5bPCZOqJ9vb9KS6E4oNYnzZkb5OrnbFLZ4o8+21lI6d8tx
hT39XAYv0BTLAALRpVA2LCuhdEYMc7V9nmTqmsYLxpkFUjZasV3M28yIwO5rf8dXxiDvxei4za5n
gRStKC5mbSLC0X2G1zZqt2/AWhSJOKALATrLb+MYbewdVfRbOxsEReLOXJ+OwagfiNS/E1Pj/hGu
0vJ5cx0mxd/HqAGhjiOA2wQJuVcArg8i0LjHPKYbvnPUqTEHqTxrpM6vITwMgkDIUMyRk85siVyL
M+zoTkFxUa2YJCxy1za2DkPHgOXGjuQB2QIW8xGNvddLn/jj6C44a0XVioqV5zqoo5Bh09hxZgW0
zQDrJMcma1hm+OD8qkcEmDIpT+bOeZbnLbRH2prYkU59G5FlN03raPX7D9eJYslM1ic9oKwpwMSF
iaaul93oeaP4tLwZl8shoNLlLHAuRlWTAGs9cdsrEQ8tZubFWfpHJ1qEuBLuNp2fC2YIlQ3CWvXo
PTSNkWHB9/FdEVz5WL/hQKXAN2822xxU2wlzfl+6Rm59Wv4pINUdoTpSUSmZFTXU+fdtKBwwEroI
Jv/z3em1rhdk8Exdjt55wrinwQkoeiYhVTYo++LB6IE3hII5Re1gGU/PKsspp+O+CHxeXMlzhUcc
xomkIEFi5OTFfKIcHnem1FnuGdb+WgfEVOgJCyh3zGiJb42KiKzJJQ7VLB2YU4CDPaIA1VssnwtE
vYzU+Ne2+nvq9S1RqaHKw5FgxreXHGvc1s8cuyIxeLc64eBPC17LJS5I451JqF8ZrU5ahaTK9ni+
k/0nrulLITq5ppcTD7vY8vS2U42H0bKt/9caTmXyNti/MQhtnRxedNNH0isuUDLbi4VbjihF3Lz0
NZ9LZgw6Evp79Y75rF5LV5jFzZk2Z8BAgSonXnoRzwknRPaSfJciKN80J6D6SHYWInjM627agi4w
2uLBymDgG1mXMvSmESgQc4vPCp7hlVZv0suov+oMp0v3pws6aJ6DfFDzBlLP0ZFs2oIC/YQ94kY9
XvzxKqMY6ivROOhZz77A8o/zB53U7xiMrde7Vz5N+jTkBVHEhWsL3JTY0IKKRdtZENWkR2yjcmDP
NEnM25I++jKvFqsVucEUwUyUgiYTthJwZcQCn7+eqWmKT4kWEZ9qjWZ31/LHbvVh0JI3JuA4orQj
3Oo/5HURVlz46tPriu1PrgUbCDVXz8x+nym6pawGHZp5QgNHM0n+HlWCqkQtnJtbTKp/TMi8sXYd
z+Apgv5ipvBFCinbtpMy79f+XuJ8KHBmBtGFenFw+NpiHzJEaDXEgdsmgbu0cWrmQDx9Rp9sQeMR
B4yvKCcobcmx2zHvv/SE8L5VQiEZkav/vQJop3zzCB/4hElO490WDQ0a/TRwUwbO4knOp/IEC9SL
Hnss3cb8jpeYSTzqUYsBdAm5KIS/i1+PL2tW8GP13+l9JxRwQmz97Lnasma19RfU3+1e/a7YY60/
2YsvdDUezz+K21Mm/G6N3awitm/WRs6mjI3KxpcnsSJMTkbFh1noQ8qhn/h8bTyZsk3qe72AageX
Bby8+ICbIemEQPu+eo+j4JnW+6L+MARRaBToJlOx6oCbpnshnZ9VNopIEVkAb+d9ReI+H96VwKL3
pC0oPiCBX+YX28EG1UmyrhpBl0qf8uxsptfK0+pCtU6g8uw02nwSw2ZxDBON9NHjAOtb5V+AKLYr
Q87Im8KfPsXd28gxB5Ix/fWIdRrmvbMzV7UESFe05hsdG01fFxQiSK68+aM54rV4ywsuVrAFlvuZ
XlEHd7BAVTqZHKMlzB6yHb4pp5htiuxBCG+f/ZCSccYP3OjAcIguHl9l2ERNRiCW6QpQmexFFZC1
o2BTFWyiRnkAo/GVx4NZIpgvJLz8rlosQXHKDVMRSWt0bPXoHStg4MT7bk/4u5/t9ANMd7zMikmA
4SPxdWytWNMVmzV4bXcE6evUuGtyKwE7u3VucaE5aI297y9ipWcP8wbEPBOWays0Yg7ymutz9pwY
7ru9j0Icfl3ndEPyzJ61dewODn18dn8wtHQglUjmNUxj04oyBhCvuOpffQOoa5E2Irv0AvB6s6Zn
Q4glgkLDvRtnmz+6jbmks0kLZ5wh3Ym8dhuuNuCoFlOxuCZYORg9fZiawor92U6hDlGqiP8HWeVu
KDRT4diKIFacJunU+jWtCgxBL1NOBAWYtF497Ed2YV6BJELEFPXj5zt3rszt2sWN6AuZ9o0LxwTZ
OISNr/sCmlCiPP8ouolTFwf9Bnr5x6BC59pBDnPjWxwLfBHrbMWCVr0hcqKFV2pveUJluVvfb1hc
5hJugUSCZ0OgZh/hVSspmEjxbLC2zT16hk1fDooW7rvpmwMKqqDCwCeqUxn65vjdoiW9H5ukPlmA
FxN/Afn7azhTXC2r+nOYGLe1c38GOlO+/zy3NKHXenwwLTeBwnZCGx0o7AFmN05fVzMt08IQasoI
JvBU0FSiNo9jENzZLoX/WarGXGnXh8tIzG2welSHfbfeBz1xYLiKmxgj5XDVPNCQ5Wu4mexPr2al
urxSiqpbNQi6AXrLEqoO+5T/SjnEsOkZU4kfe20bnFJrFJSo5zQtRhCGUNXiaoPzLt630ZF7Kog+
TsZMXNQpgU8bozhQfhdhQ5TW1lrZoFsG6LwWrC3iENp5CnDUJW5sQJ5NGyRUu6PejxE4W2rVRuEL
Guxh7+pekWziZmE6FLNz/cKxjnUJyIINPbY5e3rjtEF4mEG2XtD6ovqQZhuOBWOTs6Hk8dwH/g+M
2xtKoGgqiXybAehziU+SSMPRHO7W17wttexEFyvaxOTvgIXbNZ3ihEHw9Xt2qi4SIMKVqoCPPJ9w
UZAa4VTwkWdkqSNHVLhx0pVUV0bRJN1T1B488nBTZ9mG9xuKStu4js0x04XtFXxUi3JfG+xPl26C
FBZmlymsAgONDkkpWSLI/KO1yj5s7+oPJh1rKea2/LdaHGZTbKL434DvOsped0YdGqH8hMdDHueG
RgO+kFbnMPRLdmFOut9wdv8gXRRuOtCKoLG6Gumoyv2QoQukcl5WuhVCW8gA4XMv001qVM9rwVTD
N0HWfQplwSWhem0zMfOZQpO+LmpdKx4roIqlVW4wwyHqIthG1dbogTol3jAvl5n0pHigI9+4szEk
jZaT00p3S7RRfTXQ2N5ShYmFVxbQFwqXKYxe9kCVrmvthpiWg1muslOr3YYXGhVijgecBxHJ7NBL
/7ygyOdZIxUV/E3eARQQ7EZidSR9MjPuUsM3DRdwCk9EIFgTXb3Y+LiGrzzC8lYvUp2a5jgj+K/m
vv4durN4o6va5/GbDxz7RSnLCbocTT7k8klZduybOhOo5nGeUuiVN35pko5+f2dgW+i1h7PykqXX
s6ZV1FsrNofqamBWMYJsmIk9GXI4vtdsTSC0JJ2saCmNOlz+e4jxVtqPpMvn1QehfC9/DiL9nhrn
XrTwijtJj444ecrDjsETzeGRKLXte4xmQccSBhrg+3PenRTBYmc40pF1lckw66HSLJhr9Wsmd98r
Xcbr58qIfjFcuMCBB+hJ5Zrv/vULnggq0K4GMw4TYFncsEjGfg3giUYK/C7ilDjottw85VgB5cRn
mNszw847X/6WZKk5CpUPlQtFcTsGTorxBsePyNiCDgDM1/TEmhYA8PyoUj9UrlaqfaK9PgGu2zZG
AW5etzi/OfBZpks2+Fprh79Pi7O1a+2VavDWm45FBSzscX1/XaSulWcqRbt9aLR4djTqSCKKJewz
q2WeXeXzBi2DuYDgp1nULy5JayirF3Zb/5ZcJULQ1aIxSd7I3NAJ6fU39hF0oUX36S1wKUbGiRko
nLtY5WUC73VrD/NySExPcyMfCFg2zz8euLKFe9QEsO6fROu7hD6thDduJHr19Z/umQm9iucmnYTO
uBwjG4QQb5xZaCxbaSPQEpwmUrrsvZZb1fKykgMoEHRxrDzEkFWs3ZmrjZnNl+uYY7s1OVZfEKQN
DpHC4gbxi6CVBQFJPkx36PDuHUuQ/UVJMfdaCS4tC3mXbSWBXO+DlysfC6aeWvl7RmrHdtxSvxcp
4mdvshyUNMAgjvqg/cPuGNCIf1nxzv8GOZ3ca7e/KOmZTDF26bF3b5+dq+OQ9ohGcbFTZMomXyxe
2VDYXtJhh3jIk0VKlAY3P0y27gLndEx+gAuV4yJZkrM9DxJDZoR3cqEr11cMbj3g4QmIWTVTjbbC
pplL958TOboQqV5tCWHnhF5BSFa+t3/wsht851j4Ay8CDTSFS8ZelWGCCi2N2eYoSSU+OWWX9qD4
ozf4LDogOev2Uoi4RbdHi5PRK5crJCYGUMpFgfwyrhaRl5ia7v0DmUeDVxuw5hDiFh622BnnOn4/
JNQzZiQEdFLlG+GlcQQuE+OCr4qpqK13obN2GAlT49OTz3dyhu5bVHSPQ3nlMszIJBt8sXO6z+kD
+0xR10mmqrMsQhHwso+iGBZJ2WFacUdhhJf5EhMb7lLJeft9XhUfVAa5yq5D2xrRDUK68HZETfyd
iI9NqedpkhZiKmf6Lae6HYA+LoUxpRT3Mr89eJYcLW4WHhN/OKksWZ1rp72uevZbeOYDRoMITvbZ
44oUqn53Z3soyCQ6buP7QdIgIwG0+wsshH5nase1zV+RjiH/nuDtn0DXG3NBPdKxDE3uD8ppVxYs
yu/n1B/VciRDbH20LojZZ8/NfFtrcHwoSbLgbL8Ocu3pFjZ59uSeD0WnvyA2UeMSSYUbiUZlSsqj
WVF1PmuAfv1ZFdcZHrT9HuLOuLA+YwAcO5zGANg2/dlGcWGsHRe5KqWgSQEfb/P9aqvdUdgvd1+7
Lc2fBPWSrdjmT2lr8Gyxh93CPu2Bg3m6DaUs5ZqdCGjJZ3Hcn2J3VOkf5c1DLAaihimy3Vm4+YY7
XRyyteSvIECBWbnr15MP8RsDuDB1YXn3iMpMENOM6G9JkrfdN4Sn1oRsS1Xfp8xWDwNSFwrDq0rU
dBjf1HfbpzkDn2sLomieSAFeS8FQmkHihZ4OGVvNwtLnA4kjYztuM5mljNYz0bbJgjWsNG8tqnLJ
1ASN57hF5W5HuNZYuMF3MjIIcWs6Xx83JNxhxkohdbtc7nU0py7nuEUqdTezQqN8hUaOQBWLnkL6
OCzRsK0fKt2LInM9iTKjKY5uEIM59Wkyz2yD3z2S5XnUgDjsZ323vSY8qwL6Ph/xjurfA7rMEmxK
4TnQsCW2hlnDIgtFW0au9lMIcwmcm4LMqmfgi+x84gfjHfIibgLL6ObkOCiy9nFLvpWP35L2rXw3
0khRgfx5SfMsMW6bzqTf5MtIebXdBFKCJIhV1VGBJEpYXC5MEOQ33xoKDvn022i2RncdT2Qy/CQ7
ZiKfN7kKZ6wkk/PQtAWRP1s+lMRdgyEZAjYTgSScismAT13GDNJe98K3m4GY5KimIuN1AO6oV0eu
2EIpF2WR0WD8a0vxS5j0rFoKJyMNfeDPCLJ3/2hussqzYVrMLR5pOIBXIKOxu4XlQ53cU+4h4jV9
CJVSf31jyykh5F24fj8qONqUrUmElgYWhEzC85w58osTQgOJQUHzMkNSrQs45efWQpjDeqyugzqL
bkYqKZAcJuIrE+rpXbcwsoaVC81I9wt+ocFoTnxczYKlfZriQBdXrC1yufUip/zG9BY6H2KvhmE9
lYLPBgNJSCaNrkdzRPPO0e0pcQST4Hq0510+dwyjMU8W6r3Cw1uWb9Tw1QU63NNo+yVTFg93d68y
wZDEukqwqdpmlfFxWqf/bAIiHAD2pbdww1bM3XMEIIp0sXZHnJB3COHtgCxahT4KeRs6awGAq2GA
/YnjHRbFFEIhIOi8+VjrJs3/w0sf+0y1YvcTMj8tWmIJ8DgpoZUpZrcGq1fMVHv7oGRkzz993uCT
zeeO5VRq2htPc6LZQaC9Ap2G6VQOBo+Y5OOoQe9bqB1ZgI27xIQX51ZpNeqA6IuM5lKnJon1Jv3i
TPqqPXuxmgy+69Ug2lMWYe0Z2v1stRiXAn2mhP4a+sKkc0DNyS+TdU6rgcHsS8vriHt4Z5CCTESF
ucz0siEH5vQkgWKeAhBa98KTghMt3UIZGYM3I8Exf1qKnQZfiRu+C5lAAX1dSngd2mE9EHjk8Znz
ToMUWlXFstGs6gjmEb54Qwm9rYwQsferYtXl8LOHRm0vBGqE/h4y6cbm0J4YqIQ0P77IhXz3akoK
OxZaMB2dIOrtKSy1a2vffTt+d/+KPVKrH10OqCFK9m2przalx44nqrLGEejmNR7znl79yV4RGYpt
87ksefE53jp1gmIZtzFPOJOnJoaCwm6mCeK0Nw/B00cbmwZFtARURCqgz94mcLTy5CvrWnRS0aUi
hbTr1IrRbtHG6CedU3WJ6P7s9bbEBen2j7/6k/YmAdoF9s+ZrjnLMTLTL6RmemLNoihT/wLR9s+3
oJAbup3wm5jrF3fNAiSohloC9aFDn+kTHowZvrp9l/ZWlfCPYVs7pcCaMaUdnumo2XD8cjhYTAoC
Y3UdOkzHgqXPNhQjA5wvlalC3izKaQQ3OBPWpQoWil79Lg7gITZaou91JXI9i9UFw58+upYGrlvG
Ezp7y9cftDkxG94ns4VXFM6L66bqeRZbi8glzdU/XSLnpfqxgGeZVNbo2lqtrzkGhgRiFsVXcyUm
Jdd5poBAV1ybM+BJsUbU2XOTdrueP4geyeadw3KNB8phx2Fn7C348oO84/X2UYi5hfNOOJ1ATSDt
Vt0Kx0SLWXMVn2oV45k+DjZLKLnWW3dqyAGg8KgKD+pp8SDh1Go2mWCsONAv7FMPjVen7lzKQ3lp
wuiuL6c/kyRPAIwQaJL9/lGBDzuXN4dKSdOFeRu2GHm7SgntHk3/DX6PrCTe4HS4Q0QOcJuiy+jp
eL+MFiTGEu3dnwLBebpv4t3ijelvVxKFER5yLls9DsljUiF9P81Y/2ZMNvan5TWFKYdoD24TSzE7
CGKFNJiJKQkGqQCiEtD1hbssIJsb0eex61wlsa/t71Xxrci69Ma5sr4UKQwsAfF9Qh+UD+fbOiW0
oTXO8K7uhcUFqHfsvLhWlXPNgfl64WKNda9Qu9/iZ2cjEmWPju05VH8xYDyMGZ6ahGkFMT6P0gMZ
lfaxZxwCSpdPSlaC+qnCxicV5U0TPdUDjf+zMFgD2R6voo7xad2bYJ0msqkRE7vWEQprPUcou1nf
EnPvAKpHvMtd6fpyMZZ5DesK7yNPbFyVUxkaO356DKT2lVARG/9AlRxR0OztT0a1nSvbqpfLEB3K
AlisU/DW/jOqdj/KrAFHgGbqYVvwafbXX9AGlawmE5ju7xBt6JNYWlJ4JGNmEJkIKi8byIgRf5j9
tRHkKxYua1eRYyCOI65NsLPSKXXzWlygwTL7R7MOrQvrc8zTzsad1LnBEHpO3W0wnOz/OSg6WEu5
ITKYM1RtYcceOxzQ82EoBrq/bTCqm8UryIWxZXjBnY9mHoMh2Ef/r19UBgdmYJ6qxaiBveP3g5ua
oCiNDlRmoy4BjlVo6RNQOQpRHXGhznfouyYTROONP1qd5FRS+YjbIsr0uRjLPmQfi8NqkzyN6QGe
xT74y01W/P40DHUOPRXemBhq60hijrhl6lRrjM0gzxXUKaID3eDJ0IuxJHcbtaXJioDPuFGprL/L
9LaqHzPR6mCWlrKCwcJV7NyJmZp3AbaEoZXAOxE29kzCDpU+YhPj4PvTYHprj7PA61BH9CaLLaGC
pa1XqUyA1XWSU6IzO2r4GtdGyBEsNDhGtAGcw6SCctM7JgdXGF/2nhGsuLj8zWdG/eVTaORvSgXY
Z8kCpfi5dpa29TkBb2RnP454CX/DA9fL0y84twdiE7FFQDiLbdr+eGgh5bYT6LeP5UF41t6iuR2k
0XC/PKAAoXTPVHqZU+KcXPUblXXdrBgN/m+EqhnJnmDISSNFIMI89MRTiDicR8xaVBSn8mJ/o/0o
m8hrDLQ2TGn/FzEDV+I8LoEjKLPMb8nYaTDhaxS3GeIrhTShUzgkvcic/mJ2XXt1ZmxlczMG8vKC
d+B8LqKjsWEnt8u5S/SXivJR4BOEIO2kAbTDQq6ioANU+WmENnXFcHNoViV1AjLorLhnmoNDgwjm
YY9Mrz2rMi7mzb+uIwEmKXdEU0Sf4yHrGyR83Cwq/bdjCnIsfrkyB8rYT5ezbUW35x5X6IuWw21f
U3CZNU/lA4hOjmnbCYO+86U7MVzIo32cbFTfAajfgJl5zmMz84EQ42WJwPLoShMFUt5Vr+vje4km
Lu5Ng9ZQ5qvCIsf4Nu3imRebfp8yOiQRFi51gSK/dwQ47G7bZumPZlTbwhnfbkH4/HSiGZ+XQb5Z
uP/qERMMi2hTUIMSTPG7c4r7gvluRQhoMxlEtQuMwSpDdkFntERcKL5Zd6MxnNJvReHU+KvLdRR+
c5vUkWpcakolatdeBGX33gK1py/yddOVpGBp19Q5lRZSpWpY4JpArmQaxfMAWkn8nrT1iTaOzaAZ
4GsOiu5yOO0csm/U49r9R4bE2sU/p27RXaxe10a6afW6/y9XHKKWkCtihAMAgIFhiWxf7Q4V3Cnn
3TD3en8d2ga0et00OTRvmySkDDOl8nQooImeVHccDd/pscRHAOMVqm35eop6C2s2RGZ6cPEpmJ7/
U5fC5OIGk3KrqnmemBXMUSwP8soX/JVBO5jIQnrIYQtYURdHbE3LLCUzwB5Fd1yc5d2MrCR5PSFF
w0ULrLfLUNEzNuIwllOqJzBd2Og2tUBmq9JPWj+jToCmppdIWMb9noo6/M/xjvQNfIrkP5lzcxXD
DG4LPeYXMLQfI8A3vNL/4KprE8vbBA7ScUMxLCV5jbwiSL0B89ltcJBVhQdX+8e1ENbB/WNe3xhZ
hLUmFD2rMrwyynDCjHlVSI4ER606wBTcgR6aP1hzRflR9Bfh86MwVdRsTWjyl4eo9zfUI6ovGGlV
KEvpNyczu50SV6R+EtIhVJZ5PyZZ0+1fRjbSCG4q0GqS9od+zt9212dgI7FZgxMtOZUA8o32TqCE
u1VbKTT83rGQOuARfKn647NL8S1KdMLhVRnDkUeWekoWEWzoPbdiv9wQ71CN6Da/V8/LR+VD2dpz
S0L4GlZfs0/zfAjD+Ih/KkaZZNkM9Dg5ff+FjkxbGkdJnlYhhuxt+zqa24J7ZdRu2InfPbDR0Os7
/r1mpJDisdS0MO/hfyDGZYkH8tUv3+DYvvNwGmo5RCi4/Du2dIaFcouHTY5pI227QWSYgd6waXtF
/4huvQKBXSjyV3ByYggENm6sr6p1s1bMtb7HuxKddgIkzq8s2itWxYRvvYNQUUObd6KMmfRodhTq
CYtpR6pFJsScn9gIIbI1O40pdlWt+apV47m5EMFfFda0PeSdx4IkvIIhoVP44XgSjtISU+fCoB5K
XfWhsQv/U5BWJjKsB6zw6lYgVKPUjYZbc3LA059Rf50drLs9Je3+XRD7aatyv4QnwJ1maBLBbyFH
HBe56ZJCgc7f0mzIYEqm8LGydrd7K0BcaH4a06NL5pYghy9Z2uV1iOO9V7CG4DX/Ab4EE71NM7hN
Gl5Kf/HiFe6Io8OObgdxE09SqP2YZZSkLnMjbSneY8+WMvN/nzsKBOnkmqmH/yfiP55ST7LxX7Xb
FSeUb7D6G1m0BKSbwdNQ85TvqXZdxuJ2DbJblhCI3e/FlG67eGJCae7DauE5Lb2SroovtggqbWMS
t53cJtcZsFyoUOcNiY9n4h2zgKIiN5L365h0KPJjUQgZrgodaOrd4MfI94eFdu2wQvagHo4OAE1L
FA11Ri+X5eu1lwJnFNbmgKJI7R3Ot5AkHpOYH96dji2pDsZFytLE/9jLNkbktu1o6gvw8m4XIDYI
OfDAxEO4KGP7dRFJsxotyiDd4FixiCy+ekOqt6YtrK7HL4lHdlWn40uZWgC4Ek60g/OvfmPnuyYp
wOxM/FJur93M768z3uPqZPjy1adDdKNqKYMnhdr/Y847h+lH06oMOczxv/ONkUs1cyji9uVGNRsL
EJNcigYWCelfG2vF3yieRKcm6algnq11pcfvNZ5HZBG8AAsNLT3LczWnMm7/MMWNvaaaJnQXcHIS
c7MLhoXxq2ZWlNiT7N3T2SF8cAD6/PNyalW8dZpbtks20TtUNwycZMq6u8Ph+MapYiKdbmZ8kkTn
pmwtvyk6NHzTdL+LCjxEuqfNMgRlWbppJ792H/5xncBvcOm1bAqpOSQ4NZ/lPq+eWd3ZsSMdmxN8
YmXeptDaKFRoQ1Uf02xOeA5+dYnxXsG9bKHtj9f1qbO5H5w1I8hk9bUw5vQuVZK4js4Z7NQ65Nwe
ZOe5XJkqs4oKyi0P67VgsVBy24sniB0qTONkeRHXgM5cwPxhFtkNNR6hxwYLcosg6bEGe3M4Ulbl
eKdWu1UulRdJ0MKWd0SIt5Ak1z0gxfUk3ta8Bhq4HbTbwGVJpOR/9OmUmuzBUXU78nDWeMOj7m+C
xONnBOSbj14jtUTqj0gK0NYiAbbMGJf19SFaUIsiWu7jkM1vrZKsCTwOSbUCdygf5B31kB02F3Hz
bRaUolwczPpDY4nDTmLheO1XBxbPmijQd1B8h30mrQHuk76+O7UE7IzAEnLChdtr0XGXumKpIEvH
nBP6tfLnMGaZFD16gYQqcnIiklyqAAGfKNYzi8mzx5NZtTnb2s3yVPhl8lXbK6ZZr7fn/1f5I6EQ
MMY0GT5KIfOYNnVDmXH4dL/YF6o8DAsSlo6TuJ85Q/fjI2nt9lgkInMQq0mK6ezAJxpdrGssJ+1o
5WEvHDNTSd4+3fjVgmNR4DJRAwM9C1eqTDXrDiDUQna0sy8c9IhwW70dguiIytJvecBENaq7mW9B
tq4d/mCToOwvpYIGpmOVN2AgRlGGg8Hzmz/HThquRZM7DS31zZ12LF/fi+EPdE3m0x3uIrmTGybI
5e6Yo1UWti0PemhmbMceWsYoSIgiXjEJAe2SCltNG/r3WQlalpE4YkV7F56JRkxLu/cQ2FZE4mqm
dfssLjiTpaGszT/a9+0ganJ2zJUeKnVnBcxt4PYBWzcAPE9Awblwm3qVdhp9vFLHTgE81909MtWQ
Jv/RRGEKr/PUbL+cA0vMRsMeUGjVI1/w5HGFExtkLO/ukomi0cHL68+01N3974KSHS+gN8BuMMGD
C01YmApvzT4QnCnA8sX4kz7Yef6NsD3dZ70Hk8ZhfEjxtnMTcxo5buMFTCFeCbDpCE59HTMSqMDX
6TWRveGRuvDGqIRNec0mqXD1wZOaWm9XKQIgUFjM4QPfxvv+WvKY82SB6yl25NU9QEIziV28aupP
HE8qqWlAA/sL/7whu3F9rrO2IP/3UG+fUrcGjTcawSuoh5I0VJdfDoh7cccCg1pXXooKgUleJchN
Ybml9wn+jNj/+uF7hmp8XRzjOQmyVmQ7+s5xvhkvIgKs380SbbixA+MFzujfgsEEcX1LUBp9GzUq
j/nDC0e5dVv7KvD2Eg4BoFBF5iu3vsvqxgIovDTSPZQDtafax9kKfzzRPoyA526GlCXSHD39WAsp
qKyQk7QsUJLwebjfOWoPfhSGPeeVUIBRM3H7Ze0/opxUtb1l4nC0EKlhkGO6bjUEnTWv9zUt5Ri9
0fwATKNTWRUIEmCkr1w7p/LK6bD1zCGhb6TrefzixTOrzaYRo7L17efvzUXS14T51J2kudkPGo4e
kX9/erBVh67GSOBUWka8DQYDvsL5imSIrgMBD+lJz2o4EvyYvmRrXDaEkObhLVVzlyWeyi199Ndx
tcYbBpPLn0KZA4+zU4884MiaAQUmnE7R+X5vjcytDHEcFk9JZPm/GgxhrCCa0QLxqHrTh1+dBBvI
dooUY8JxIn35bYAuQrX6XP+Q0PdYyLk7vC8geDcRBqjnQZLVDhYYVuZKkHr5yn5DG75tEf9yn+w4
cse6E0JbUBaNgNuHXQ3I5LVrpqORjlvOgJq4rCbQE87DkCXE/0nNoVnP8wS9GEcQ/OeJS2hkW9i3
QBTKvxQIAoXB5UcNotQToYmzHA3vKyfmIKVvLoD4s2CVqzJjyH7Yjl2usqa0YFP2XeNON3SYMGQK
iW41vQmHr+BxZFql7G7Rhgnicx2LcETWMMhVyHw3PVvBN3sCaIinxBLOuWK6jowuY5uZCexcA3PQ
ZB+gwzAghaapbwCh/7QGl9UAOd8uNLoo6dWRrRPt8tcG+FQRaxNIfVtA5NbmcetfbRzjjOe/dYb0
xbq5g41JEI51XvBFEb5VcW2ZHIz0KK7vXdb24Lrjv/qp+RqR+VF+lpfqYZmgRkDeWMdL1f9J1wxm
5zSXkU+jxM3LBZlR869mpQFX1C2LgZR+ZQtEAdUtgtT7tmMucFh15VkmlltG5LvWLY+KTSMNaljy
3VN9OiVrNE5F+piaCVoD48qU+qLdDdKGbCtcJgAtsRXfbi74P1tcPpxjLDk62ZIvpygfQDcd2a1q
vfF4/bUIT8NjgKwk0Ht4KGnBBEWPs97x14qfanBflkn+vW4e2faL/zzikbSiMiJj8qFKrgJVFRc1
5oLLrVWH9CYgfTLG8p0BAwtfhXosRu5h+k72phQq9/PSqnhdGxFbVQg79kz3ByCV2sZRnLot2S2X
iW2999BdDLQU3x9uyP9KOPbKTUeHDKnKp/BEIaH3zl/a3c7nBxCrfdfOrz0YWW+wAxszqvyey2go
RleM4s4oMy4RPWUshYyuKGpO8KTG8cdxmV49PDD6wMkwranmzvpu2EQ7N70ACkpZWKIP1rIqi7wT
w9eWqoHLu1kxxw/tjEuakkDlnfVwYtgTppyvtHAxw0BZ6G1Z9kggQ8yo38hRrVR2IdA7JQ200cer
ALV+MBVxDyMRVDSyYDM+wgNM44eT46eb77ZlTQm0cJ44FU3v+gO6HmAmnTihvl8YqzD3t9B1A68J
i3nCD2ZDbE/AvVplQ6uJAov1K0+bhoA0oNx2eMmg6ARcw6eRVe5d8bEv6PQLaCFAcoIgNGvQouwI
XvutBA7155s8b3SVG+X41rB+TupsGuw6LwB1rZCkBWCC+dYb1jmAHzZNCKYzMGhhLes4ZpE+eFij
sIxcixf0l8bNgU20FrQi09AcLimBN4XAE7yMejloVlDe0yAxNAZDGjboPvnCJb4YwMFlktWXFoza
bBCvNR3ycVnOCp4nVfO6FBuTgVeOHfSvHXmy0zVmVMmhZasCvp8rz5Fc9Meo/co1ymKxqQFGOFvz
6d6seCA2HUVFb1lyys2Rvh1y6Uc7FDYJEwiOCK2KL3F5dG3uRMY4Pt1M2dPqGXiAUaO7c8/Tm/y9
3tC9sbksBTVJwXIqUyLdwoZuS6DEXrc0UTu2piXPBmdBxjStmivrIT+RzVGCJNlEaHup95CxYOHl
OdepBVlr/wI6I1QujqSUs9a0axpZVnZZY6xe+c3vU+BgiyDcUPFdwGmi3ni8Y3KUsBxmP/CjaJBK
/VW6LreHonMvjzAh0jFAe87ujT6s/g4WvY29RkjtRgwk7VdVIAfs/dMMS8XOf/YC2kZYb4BfiQlJ
ZGO0TMR2n4DXoGdGhy+z+z+3cEBamB25FFF9Krt3fY7FMSk9B9n2xFxac4jrQWrfmQT6Fa/HGssd
2ZmRNNpqmA7hejdpEGVmBlUL2XtAlX4cwEn1Fy5aF2xX9KELBg/3hpgOgOVS2YSgRiW0U/Sw5dBN
aKxNgVxBiWBMPP3ZzMQ4Iw6mDm9aeLr5m97OszBtfcinJAOu+0pW/3pJtMFpznrq8j2ozuSjP9+9
TicD8e4T0KJ/ZaLaahQnj0Hg9rlbV9uayD43KjwNUVWnDOwL/GliBNm9EtKTqQTRLJ64GoQQA7J1
JpsqYPoB2w2nwucEnleGAVjAUWV/FS/YsY3EHb9m95KvpiNYTpLNv89skIgrg8ualXKnw46poFKP
1yU9GsC+p2NYRrA7bNxi5QlamJTAygl9xm1Sx3sUaPrBgfzqgh0q3AD02p6msu5BOdpfsI4uykFI
4RDyxlQY7PVDYibge5ahBqQ8miJOqO/qJcp6HepPkV2STTB6OoAf0xJFJ4p8hvnQYoJeMlXZ4Nz4
NcJHlo6CnTdY1PW+e8lLum+j1WWWzxMlYl8JsEx5Gv/pCNi1U3t0Tt2NURyuclsGXXlL70ety6P1
uu9WWQx81vBuUhL6UUu69aYijVttyjWfPjAIspkZ2NcgaKDuUBX5xXRwbreUs4H0S3wBQ0P2xwAs
2W5tibEfWfk1caeS4747n/S4mjRXOWQ2gTLZG93aU8cEvtESNC+s3ekvn9oIeHapfo3NT8cigY2Q
lc4qPoFo2LcYWF0uNDm6ETWLuANnEXVuSGwZ6Y0R1vdgTvENFl52XXXTlYZpkXTAaVQFHZ7mAECd
cRWhjLvPYwwxdsJzS6eEl2TLZcwYVR67oHRJaBdzZ5r9QEQFPXTg+8Gprss97Zfbgq8kviNuNoMb
42T0yscN715g/Mhzgd3rwccxiG90aMNjE3jU8s/mW+SrZptNqKZZwDRwcwZWFa0hsg/05iKWwNJV
rWm9S0zzxMCn6i2iAcLt/DGSZVwzep1ytm7lvLsuN7nzDktKpQ0jmjUW2aqvSwjsZvpB75ymyY6n
BaaGLDvLJji68Rc+qvMj8nPXH3zegfF67L2TrkQZgJ4pkPJ193DpyXp5S/WGyM9EqPuwKivulCr3
6m+wYkwE1Pt251FbwBTYkt8gspWItyBpN8nCEloDwulTLMJcPznaBJkPwgB8gpceMe66FnHTQ4yn
lJO4j+PAjGSh5f0RQFg4rwztavP8paUfZDCI3t1NwfE3p8S6TWplQKbylMLTj8088RhVJdtI9mNG
hGcXcLoN1o2hrTq2R1mfd0AKZtTpZGV3b+UAU2GziW+AIbS8NgmE726CBFXK3BMv1ywdkWLYN2EE
NhrkwXnAAKVYnIVWcFczRDq8/66PUiu/2AnCPLHi3VgIYNl+Q3PYG06DAAMHE+WAVrjyahUd6Odm
zxYc7z4ouzg/f75LY6tmcntdI/IDLesjXQ3x6QMr3I1qDa5jFmbGfRHqNunax6P41uO1Vu5Wwnv1
MRzmkvj+yo8XMFZFmNY+O2nb4NLMTGZ+k8PSQpIYqS9j7ktLQZsOTeGHH10xZYyUOmJb079XkMNB
C/9mBrWKV4y31kRJj+p2OzT+xYM78IkrE4UaIT55IdsEMVZH1GPtK2GH2LB+ZtLs4ro7ucBCn00Q
nwELAAgdFLrY19uHmdC/W9Zx8CwxcPCGsgk5Ore9YUozxxUY4AFD9lJP/MCBXTY7OEWmUq4Y1NRA
aYSSlQlbg8HBuzsOaeHhVD8pw2QNwWAKOUG4SW4dOl497LtUlaAimdMKK8cIUgu2UzuNsrj06BEY
t13gXkqtoHeh0jPSbLGlX5thXPE/AaAU9uwPzSYzK7aabhCh0EIyakwU4j5PAQ0WVUTTUjMmdKgU
OQr13GNsiCNQiiNijm0zRP9jSl7cIx+zCPc9r2REjmXybpH3OmgV0d6iWSS3q5zUnvLrXB4MsAFn
gAOmKZHjdFQb1cUAIpIOk2hHylpW9dm2LFrkFExDXE0vv+aaf7KA+ApNItGrR+ImGHhOdXg9oHYe
a/WAZDDW+gJDlYpPEbdASK35g8+8efgsZhbvy0iPaCtJlfLgGwyfJgUzMqZa/lzdAotLQDYd+6Bq
zGTV0nyF1LqD60MoKW3MGimjZzjEdtaI+DdsSsK3kqK1syE3Bl9CuhegGaLYklzvGMsEgR365TqY
DXiwM8s/CdmS7kx5gF1DtEOip6/W11XQ3aWQwih/3xrQnVbJnDoZ52pExRpstIN/DlwG/FrGcaX0
0IT4D7FcViGPWe9EXNgW1zNm/ojDx+cwFt4bZliuwdnid/ULs4oZXNTNUoW2gyR75IhJN7cNWQ/A
DNHzXrCftLVA5qbLFNggqLjD+Dhm5FIWj1OwJr+GCfCIuwvpM/ETZF5w8SL/71JMS6xJPBukbcxi
nN95cTid4nsr0EPQyOfKpiFPZGjrqlJn447B6GbocaM/Quy0qYabwvbTRO73zfoUXQmM9ybueqHY
MFzkupKxFIpeV9wQmKjiSpMY6If9okJgY964MsrFC5+rWsZJPwAFIP47zzdU8eYkGS2f+z78+un1
Siz/6D6H2SD/2kfHbYZ5bSSy4bqLMsyUrZSRk7gJcAuN+dUWRFepeslsVNOVkLRjUKut0xGXkiB8
FaMtHqGSJtZZaLGNEbDnrK3Qx44G1duodmEUZDIfLvPHNHGP1qx0GfJKoj7hs5s0R7EIdA9anZTq
MR0E6u2Zgyn8VCOw9D7DliNfwYfb2+CxKEPe/H6OXouyFxiUY3q8zVOjOIwS/QVmRXrEiW1P4Gvt
jFy8/QwdzbfyoxaeDHKzVs6YOXEt3Ifu0QYObdXspDZMxs0ZVa6YBClji0QPtHcr2uIySqlX9gdv
sEANGaT5dh5f0VX74kOZqmyRKsJ1GhYvUgLZikEw0jOBm/8fOKQhs/dqOTiLnMBJQBHLPx9ULbda
0z6xWSEvuEAUChZXX94ItRms9GrwCBPKpwclQxj1e9/c4daCD+XOEs9I+sePmEO9ooSFzJzzG435
tiyvYKrM6DQvAxt1lmqmdGAWNMWuohMshdhdmbfWh/VjuoEB7rWyn07e62RU/sNdDgDmYqIITjJM
eam/mHVIdBvOAhfEsQJxi+rR6s0shlq9Dn7G8qS91IAR3MwCYFPSczetzX948MJ9KWhNiNCmhrEF
beFmLvkNqk44ohwuc5ItrniH1JWG7t+EGRGgH9ypzgMxUSACPl1UQSvqMPaljk1Hur+4r2HPPqJH
uavaOFFPd9K5ZJS6cQZH7EVMoOYvskmsTnWVODkto4F6NxI7f7jTt1RFfL7XV57ENXJIJLr9VG/e
WcNLFtMhY48cI1zsF8OGi+28AzcrabiQ3RVoOaAQG7gPFhsg5865i/Jg+pDVqd/7mf2WVpio1bpo
N+yAFlz6hIeM3qIf5qfTCdrNec/X4KEUpkiYizsOCMrtOLTqcmeZ23uBZd+GHOXxpujaH3BGLN9m
9Qi6ERzlnV0kMAudrvi0YxJt4YpiPp0o1m3vFiXXIAFdxScbWhCpJ2kLMnfDGMuxQ1jQYhHFCJLX
fs75G4DDuyJo9aZ67BVP0PkWJtH74+O2up6npQledZr1YLsYZ+LgaKSsH+GLVXD9g0oZ9bgHDKK0
r1FVqMBfgZfXmYSIsynI6eYFAtcMyjOX0QvEJHkV7ubX0x6IRnyDTz+hKjj4zQVXOpshXM/jgtRo
/gjuWaa/fAiuL3uvpBHkXesuc6Jr2mCtT/LBNbddhvNcBjX2az7VLN00wl9haNppSpxSMgbJReSE
dFR4FgnIwGLUQUx0zv9fx/3FjeYtjdzw1LFWML17Zw+pnW5X6wZI2toodoP4L9vyAPxa2Lf6uEAa
E+5IzIrRSYDdSDqfOdK5bgTL5CQ60o5/qDGLDkZjTkKQmDk1oi2ZMZM9yeRSV6FL6eaA3r+AjEFF
zwzlP6ifaJAVJTT8S+erhCbYfVC5wHM0kKCP1hjBwKc3+i+9CK77yIRpjZJRiI76onqFl1N7KeBR
kTTWq0ZLVHdPMi06UzYGZvuueUuP9jrMEZKQevQsBeyrdWeQoxqvPS+o0ocyvy88jdB/LlLqTZ96
WipRTDjUKlWryUSkaSu8Jl+OnVEkb7vZGi0kbTj0lJbXzoT/3t4tjZOm/rjPJ3uDqGJa/oKkR8qz
wM3UYe0sktniQc0rzcW7Wsz/mB4zCPH89DLHhp1gz2+C8414D0ASMnmeVb7/cYAiinmPa7GTOwhU
RKZckVeWqBN3NRwHf5aGoZM6BlRblYHfQ2sjYGnh/EXSkoucYNnKz4sBG/UUSLX3L9YCbYwgB5qv
Kat6kYs89z3jN8xcDwWao+kHtzi/Oyimz0x+z2j6GT82WQKbzq2QrLkDRzfdDiMQpQm88pzjxntL
MLmAMzCK+aUC1mPYAj0R6R89qnYSh5g8D1fLqLw0w0EMSDep2yroWhwbX8T94aj33sxLckY2AJUy
q7VuycosTCBfABjHQzw0rv3KabnLueDrWyt/7C1jP2toYId9u1gGs4lfGvsQFdJBKHq10OVUml3k
xhc6q0Bpz+yA5NCB70/a+f7peYW5/Sl0xGxqJlVW4M8Ds+YoOlve7gHJa5K65AzgGdvDNDtKsrXD
UybxtDEVbSl9wdoL5TBdZJEMpbjwe/n1iYq4M1GE4wsfb3qrrTL0dwS5PDjs4TTpfUE0bc0QPc6z
Uwj9w2JNSeryk3HLI8YjWrW/VFbvY6WwJOQPkzuPgmE4U5MI4euumYr6WaSSz5u0Ggty9ltx9KzD
2WFtw8l0gIsqwZiVGNTyhS7GqsBbCT7cBdW7tCtgpZDwhdtl1j3GzjXd3ePVILG+KjugoIFsDmn3
Gg1FpILbu1fNW42AWtWDjLWOIyCiZFihxFSkqpUV2tAJ59cJGd/6eiwMsAMir99HJU9dNJ5rIlU3
yxtXhC8VlmgKcqsnG/7PDMNA56zhscJr8Ia8hFjRbrvWf4bTsMLGJpB81kQeYQd01+nMbFYIxT1m
DkPOLc20/13DtiqOuu1Md9Cs+u1wAEsaGfckggd0cfy35SB1lP61QzBzxegeCzWQV6M1FlSSXaiw
j82Fple0s5YIhsG1bUKYqIR3jLn417JipYp6iNYB8QHuQob/nRu0RWYq9SzzoeR0lggmGO19sCTF
MUcsOCHR3K+lSGzcLUJuHl2xcSHiqZmjgyVoGHhPxYoy9kGxA2KPeeltQ8jmy4I8AFUZ+XaMgdId
vHpjQMdmwokkibDopUyRKGWHbSK/l5cPpR/2h2k4HSqK5+vcVr8RJ69AXzHxxQAo3AXV1EJfF+iU
Blm9y/Kio0Ul6y1YHrGoEZS5zTt6lw/4FFo+XnpTuDpztnp9+n66v47GDjhDwLw9Wobp/vgsN9YX
42VJwjFgAtvaBJYs9etYTwXoNp21fPA6xxqbGny13omvyubb+ZQmDiyqWKwrvkiT3JJpOCYdbK6O
+iMW42FY+mHr5SNRhQIywZo89WjBJv5BXdxzq3FtIvFt7A2s9crf86hAK5cNhg03/h0BAOT8j1IX
9JDwz4hExLWXraDD7Dx0cFt6PNjyn/Y3NW5cDGB1riyjidNMaaEeQnSDIkFuGO9+3r1FFqSndSFP
MLzaiSDnVwXnWxSydS00Cj4qb5uWJRhbJhgnx1+iQtVKX17Le3ftS3hpSUPVayIVnj36ptv2n1ZX
8Qt/wTVbINPdX5B0pzYbYmDwuLrLDLPDUK1qSDaflX74itXosfGt17kJxftnlxX7W7zSaGw5d4Ys
M2rHGinNdZsUF+/o1zlyyj2+MNgVASgkwGlPcD2KD/cpCjFQFCzsOH13CYklP1vxCQrYFIRqL8ud
n+kwkT/9+90X0ZjywC13aEi/z9r9T0JySB0rf/7UOeKbat8dUba+VUrsSdWS5+WO0WTmh0xaistC
We+R9vAHK5HOz3ZM0L4xGhy70jp+GgemTpxXgShXwVDMuGDupowlcdxx+U2r3P2QlJX4Ty3LAdWb
sPvLj8YQMyuWyRV0fQV/ZMT03kgmlm1uU50CpCDy/1c3dp3RqP+5uWuLKf3jzQEBcpOkxwX7y7kS
h8L6YWmZEZdRU+cc6wzcZ315QCtA7RFiuSPOdauSJNukHcB0l0ZorDSmKnMRiZc3OgN7glMeMVCt
m3rzQfitZ4p3GLJ6+mwpGlWwSunigL0uYzW2PH4ou70DlfG8fFnskcd8B2x6zH7Pki4iun11ZzRx
HAv+GyQxJJuxnR+szY7BknJYDcatI09ybyLzNlPZlVmmKTZcfoK3asq1uN9MUYD0WnEUU/LyjXKi
zlSF+B7JhWRaVw4qmNIkIt/5E+ao1qIVy7BDHZpZM09lswS/gYe3bD/PEERnNpHCPtZ69RMZpkc7
UC8wnUY4ia4CP0Khj1o/F6USbRuwaKwLjyd3eZ9yw+sZO2VN+8hp1WlbmUhBz1sIqjToJYa1Toti
x5k5Kz3sXupGtQbEzRONBLpgP/yiKd71zCSBLx+0tT6v90Fh5HskBHQRRt1QSYu8fWFAwSDN3ZrU
fgSCmRdGrDabFLL68jHBSRhoIAqU9F2CD4NF3L9eU3CRXovRVFqeSS0IAJpdStwx6cCfRnGR3C3v
Bwt1nniNE1hDwsRlub29mCddo4YG/ApinrbhIyXMWxn+Lr7XL89keyeoeyD/Y4CoA68iWBm8Th3/
o1NrC3r2IMXNXjplSByyCATFeBEvP8/rix1WQwa0zhqphaTmlTiZXZRXXnLHgnPVRJ+ebjZwzAf0
2HLXo1WhIv6C0CrUbP6k/v6PQ/8W5EKFVRQ+YT4wrNjcNmOe5NZ2a5dK/l5Nk7wCv5TKQZoBwD+A
cUT/LbKHaNV0nUewSgssHq5e1T/ZSyo8M2wzApwKKZqd4bn5EFfwoOuPA4KvCJ2H8HgzKqf2WdS0
DXyc3TdPFKj7ubcMluwbAjNgR9kGeBO5aGMBk0w3gk6V5rhtge5kD7W3QtLOx7WDML2cINQ89pIm
6N01+zvsYziXuRTnl1ptL9M5tSIls+5aLQIZqSs7T46J6ZjgD5ITPovTNoWOYYEypOsvL5+9FLq9
KOBVVpcLgFWEfOR4kLfI1UXVdhTjMhdOb4loKpLEkOTCuy+RtS37ijLhlwozkaGrgln2Ou5eZaEe
7l7zE10q2P6TfrtJnD77zaBrpWd8Osscu4h6gWvksJ6aGC/Buq1DycuHFnnwXBvw++8p/bJjlZC5
JleV34auQ3YTyMyuugU9ZCA163YQMcqEI+RNx21t/pQn3UJoRXZHOkGPeFo1N0NXSofXIT+odfOz
oU9jMjVNXKq+i79hPRSMQUlUlDw5qJzItlVgwfwhy4feBOigtqWiiVViyuil5g4IfiKVIc8SKEHR
6XeUN2iO2ep2NB157wgWlI7PZZvNLLdK3lbInjDE4zflcXaxv0WJwe7z1ztCrXjr3T+c0KF0LhHH
1eU4SRfmCg4ku+P1JeSY1zWbJChijPXjZ1lGdojK3HbvqQ9e6nIp3kBsDlZo0IEx5OjnOQ9xquj+
AX0BFFD5ClfAMIHe7RjsXuXNnTjaHoENBvUcD5olEe/bp1fVXJI6H4yiDWaa+v3IFspD/5CZGBV5
fva3AHVXFWPHJ9sd+RyNzvCDWq82VnGu5zF2+R819R5Mwyf/E8VZI9qRqaD3yljtp+JRFlEa1RJa
g/crRDP4Vys1d+rfCFzZZywdgTUpm5zxgM6MjOzObg1IlLuuRl99/pje4vjB8A7jyPqOBMG47deN
Jr+CqcnEpCW/vI4yEt9S+qqM47OcnyYk3giR0S/Ul8yWnqpqIZOBIZ0N6j2k9M8iX1aHhqmG1IGA
s7EQ2B+TQXJzg+9iMgdbKBj9U3QZff2HbCjsFheVdfqft8tySrM1yhjnFQayA7xEjRWxbUfA8nuf
S449RYrHBiPM9O1/ZuRvRXrLKsiyhXv2O0IGGENSbSHccdmZ4AXLhOr98fBwEpmXTucp+fbhQAgC
CsmXpxvnVFEZH6kjqoVBAWxk1E7tEj6QVZgcMzzqHSB+tCkx2Kx69r9JxDwzhaMJS5mG0Ja7FOgV
LD/R33ytj7HIdiKkjKkisslq9pdM4PNLskmYmZAde+PpS7rMCnD+nz+i7XyPIPLh0S3g9xN34l6X
4Ozd90DLQ696iXC+LM0z1qBO1+nRbh2hLYEiUnk9d5QO6Sso+STp/30PMOpPvKTlARUT0hj1GTLS
3Y2LNtNvZ+H09VI0LZIJWgmKcDmxjXr8GgpvDyOs6QcbNyCltJ6HnDtl2FJpFsGmiLcj1XN7NgVc
Bm9yGRJ4Pk4VH39O6HlBZJ/a2//mIC1PjXeR7wKPuW1JzvPWVRAGObLAy2r/1ix7XHgHEvIy2VSA
u+OuvITTvqlcVXJRj1khukqjmBMS5AJa2zUeXbvgPvzpLHbygLw0DYEg0+r/yr/X3ksAtayUXB/3
CS0WkKGmDaYbLtgxgLUpnY9cLJibQOrt5RLPQ+OZdlubZ8eAy06lXeaRqAermGDZGkJskgVbrZJU
aMhkreIsxhxlOsM4SF3ZdV5s5snQBKChYvn++wD4M2HlDL6n7B55ikSrVu4s+Ks0PW2aQdUD/q0M
WVaugXGuZOGP4d0Uk7fJ0iLtlQgNAg0dOdwGuDMaHfncHfUYi/nNwayso+c+47R3ZufqCIvzMqr4
Jsg0gq8uhot99N4TpEv2qBMNuGiMVMKVAzseBc9dElQhcYqhXvw93au8BfuHzzSCf2Bo75Q6gnF8
Vs7+56MR3H+oT14zQE4E+5NVCZ0c6deO/471nSbvUXB0xuEiP/QtGLjulmoKEpaDbVbMyTH+q5vP
9BHBc6dPaBQEsUFcBOp0IAYHKIafinIxxMBnjD7GmHcgMmtOKUNGXXindEucQxmIXr0kXIofH/ED
a52fJJ9TAlZ8ezpsrabAiLERCNJN+eMIcfET9na7ZTC5FWESZYVd9y8a2DhjmlgjtviuVC1VJTir
+7asmGnr6wGFBjF6l7OI097KyL8ffkFPiBia5zPzO6AwM8fxeavb2LENYUQOeGK1JK+2SrPYH4jV
gOgyFrvTcFFCUi6KIW5MBbUDJlNhiLdgfC7kFSm4TqvddyI56XB7vrdb/XLbLfEccLc1kklLXknE
sfavgN/Lb44KoX76I5Y+aZo+w8mkbPWiPYnrkiCFG/Gth/WwS1mjzbAAVdUEg7rYLdaWwWGPfd+Q
rINrgy34HwavjbN1S4OFrEt3pujF9MOpJ07bmiUYmflzPrZjfWJSFJDZbzWQyXm5gMj0FoLORkIn
0UgQWss1LM489rugM6OIy7qs4dJ4gwrs19qFpzYpr4g3UYDBxta1PZ7WkjG6NARvjK1dPZ4X80ub
+c5Q1K6FJK9eh41qlurRnRWhb437vqrL9HKLG+ZL/s/8NEzJeLLAeY5iXVnfpIRQuLIgaXwxytBY
2ExKTeFzjRJThm9PN6L9TCaMNqAZmY5C8B7TSPEMxeKUqqAfCcoulkyVX4WNh94q5eoOrO0FtzOB
snKj7U2LTmKsnncT2Q1el83uJP9ub1i8vWAbMedISrHtMnhy8rQI2Mi3H3F6SL4iDYxjL0rgcP23
4KYaQ1wcO9Y6uK2+8J1hDif1b3zlDQOL4wRah0Ybn/YZfWLwth4nFH2FPat/uKWMW80y7plbWvfI
O+MLNIlf+moIX04t+KbRW5kL/faoZcVv5PPOoSMxjgDk1ghaWRYUCexHWoGJUhnAZfe/zU8XWkhC
uUIHc6WaHPRSjH+h7oU7h2al8fdKi55pw2Q7dO47nUTn8hXAFfhkMRlGRRYBpDLtt2sJ+TIvkdbN
HA8lRv7dhoRcLH/HGehdJHTaeu+V4TNpEUiiPD09kyqrrVJL1j7rh8UzNydCHVw5Q8wlAB0LOr1P
fJODx/enjVpOGJkdAguV7ZJzKw7ZdRAd/zxah5ppjeratrpTGxzM05PKDbdKk5CkTVUFp985WAdo
nztZULVWBmS8zNl4ZfcR5dQGWE5gXgGBvBzTT5S0v+oS4NXI0TdeoRhyxqFOJtgGo2lg3GMAnRMO
lH/Op3HTmHy0OensGFulOzJXpEuMZlFcEO+ePSGrU2sATaE8/lS4HMR7vRgfF90mjD4k5ifS+MUF
w+ttIlAlAGvmRVIsKc/6TOyl5lOA3R/7V1plo0cUxF2vKAnIEuyV/+gXn00H+gTFBsot1/SPXI2O
GpaqMi9kG8B/BChcA6SoxGWfsgw0OLcKQGCmrAdmWpEx+0TSXPcm0ZPjIwoD8Iqw2JPkv0Os+yPR
UzdX303xYjRiOVrEbH/O26ueNYuOBxe/u2mDGcFOTo6nd5rdxlh/jI2BhyBHBQrM9tTg/MHN5QE/
XdK714xF//zRji2tqenjeoAPHgEO3tmcfY0QgSZFROZcHhrReayLXCkh241NpDKALs3KEKp034cz
jUBsWIMGzMPVivt0F/HkzMetUEjErRZl55dxgglv3wQp+Q+m7RzvTx1ZZ0pBcs06Z/Th4or3z9Gc
e6MTChAgDePfbvx2Jm4Gp8U6nOjivTsqXpWjOdQWFoFg0hFKNJ7Ptctup45v+/oItZJ0+wqw/5Uq
hrVE/rEUDkZF86kewmEnL+FVH/HP+KFwFwuio9ig6tUbNA+wRap9SXVz2AUrOoITPTS2TxQcLWC9
I1fa4uqeWSqxHFDjkelPWlT3z7WvcVOwTyaECaAE23Ed9L8eMY+hpU7kcvADbSad5D7Z8FCIxKm9
gttKfDfTyVswnS4YLTLz4S+YtTvgVN/bxkpwaxAkMbny3LsXHoTHRRAPH+kU0eey7yx6hHGE3Clq
gJhtF4N9mFIZLLINiwp3yx1zobCg4tyyFlhXcvih2tgVnTOWK6MRw8TX+dBVSJ6O5QgCtWtc7MRA
sXk0Plz+Vl7tvJzhTAFC3/9JitvivQyFR7ZBZx0toG1xHfSlXKBCujO98BIpABvQ+6YAudwr84qM
r5/gKTZBDMdIS48REBmvSsaz45KxY2+78Dz989OylMnlQY7o+42OLrEWQSue0x6j066o3BanrQ5B
TDUG4NiS0kGPQNbeOJtbESWuFTkWT7GTWY8tIJCLe5PTGt8O8IBijO3gjOCb9vH+5NzcOWRnnq3w
CULa3tYOE6wJbUx26D2TNtoxP1jyaBexLPmPXam54pJ6tCTot+P0DOtD7N34TuL1Rt9q5OdFt3kQ
9Zi0IoqEQREGlbaFO4nv8b/noiyrZVzanrcW8/NIGtN3sz3dzLz6s9CshrKiC0ubjxJ06wteIQtU
Jw4yRhSfcKQdJbh/jak7l+f0q8QhFeLWBl4fNfCR9ljPLp87u5bvCpeUb1n/6lt1sZmEa6H3UAYg
A8HmIMfZ/tmZsleHYpEdWyQhBnm66nDzvZ4e5zELgycBI8cko9rIU57f8BzKHCNB/mTfWoxFWamY
Eut3jq88SU9eQKUQEn8IIMbArbSXXLV8k174uLUexiJ5wOxnQCt99TpP/PedqpNBElzEcLanG36J
b2wyKy/VOytP/rLkaDDwkHpw2UwZsaLX/nIAeDWCZMHg4QhcitVZvops8MmikFRZjTL1fGNvHcv7
/TUHHQbI3IVOgiwQAEJUOtAsnM45qOuTZ/hn67Pipo01EEfYFxA9mCGvYbnBSpCnFsQ9BibbfJ62
yE4v3fjWME81w1sCQeNiwZ7GvjqTNYKgwqdSi5tRuigno++E85vNx3uvgTsCwbcz1/ZJfd9hg/QW
ajqqfsByS97pLk2mC2kVK+iEx/bjnTBrvO/52xDgVvPqmIdTV9tVvyG9j/q0gL0s4WwJQuctjnZb
HYQPQeaRoVhTJm0FXQbTKbHNtvAnOVEtWS+G5Dv6cbLyWPYxJxXCBB9hm0x1wGUyI9xWsogLJq6J
iNZjJObGOpMUzxaBGMTK5onPT/jJA4ckdrUqXf5scam6Fyzg45wwkEIKWqNT/+ui8YtKfcU6M3co
1dto+MgqYfnvl9Z69WYg+xvt8D+jb0gwz6ZZyxevKJyNzBWrFkzPp7i3iSkJWpd/CYvuPNdEwQzN
Fvacg9YpbbVTziN3GgCp4xCxfVNd7jC56QTwGZLfmgg3NeODXLTxSQBTsPaT6rcA61PS6MCjHacx
2C0bgpwf9csxSomBK5fpF50MJbfuBkUoeEwVI6f0sO3pYS4LdWh+ekbeGKXg2havqSCeqRaZmM3v
LgWvUShrInefOJBj3EXlBRu4fzImDn8UfP0uTDhORIvQAoAV2grNvx+hGJFM8O8UOLz5qaKLFf4C
4QEk0mxtPOBTAL5N9FivdPtkNiakucW6wVZVi29vfNxvhk2xI+8zGHSWqoMrstRMIdusfGxjXBE5
dpruPjtdlytreThCJkFZAvzR1NSMEiFslBtv9m3V9+toM+8e/WaGOQCoGOK6mylP5sZAxCyoWjgN
gMUsv3rqyzWE8T0cPOTzOe16lUZBbZNfGTquZioSJoL/+uIA28hRE9hoHLH7+7+jrhZ46SJ1D6Er
ijDkRjJAshTEeWaIv0MVqPZNBqtmleqiszemEz1pIoYZdTP7dhZk6Kpxz6W6Jn46ajeKYNf6lv+u
x0cr99z/szc4iWa0seCAGFh05vynpQE86kOwj+9WnJV9y9kFNMUcgM2UuSi/rPOEVA46uEINWNcj
zte8n2oAR7Mxd/XSCjLjitu7iqTds79Z3Ebnl/kAMAybydrYikmkDL7e6Wtww87MCqxCxtGjlKwr
5ihW85pWOQzkbhAbfY5230XoLkscIHUNFi0m10V2lnRFnSd8kP8lhqrgDYJA5XdGZ334ws6fbsKW
yzUIVmWK2H7N+CsevnqfUBqsFCLsJa9dkr+ZOrOLNsRpUfcznOlV8XZPC/AHxssXs48AZYxYWpXD
HjPnyvaTfyVx6FZrUgSXTSOF3somFbZWUiBnJ8Ror8ofxsEvRS60TFF1Q4zOCQ0/Obf92J3T3XrW
XT8ZAu54Ih1nRT2+l+/u4WqkknlkOs5UhGmmSWcqtawx9EuGoxYHNKu0So5ZdXKlCHyRSMH36j7o
x/IX+n1uAz64KkyWerJhPUBUuSy1sqpBjytCyGg0SaCHhHrs5LmUDyC0XqOUdDxHnf7EBLeDLRlu
sSY764znnBfS7mM8ZYr8gzOiVKXF3Reh3UpcrMeUEqeEwb8JxC7XFKMCxOW5e6PFp15W+z2zb2Bn
umwhtnnONWOvk3DVcssMuyPBhVs7kQwUgS4+7MnAB/a9oYg5gzFJdfSFaURdqIKZNpHiu60vyciH
p1Qd/mcGwhlWcoaF+sVTMEO1L8E/0dCFZAGQDSe9+Tqjf7eoZxAeZEA3WGfV851HJCJD9N59lF3/
Lg7KCfQ/tjL9NBJrslOYNj71VkL2b16f1Q+eD3dqOwmtvR++JbjvFvnP9syq75JMOAK5IyidnxsF
Y5rsCUvj14u4ihEjFwyNTO3cNbp0Tt7YjWXj+VZYEYw9inMoy8WIigWgllfTeTnxYzuA/vLnycW+
rj2+ogkp2Ibxb4gveeiB6/A2E016vXhA5M5E324W0jANv/QgwQjIAt+9+c9sRHKach/NSCA8gISU
Vg6nmbDwLF0jNRqfEUd3zgOwS4VtDxEf+blBgUO36OGCkYEFelGXMO+skbpAZR9wUBIB9zDv76+E
3nn3qdANgEWZ1iP8IYBlp7P36WsP1OF6TI90GbUZE5NgaF0nELRq/0xwzcg4E8jKUCb3rq/NSXv+
VlCETu6Nwo1ED8RrZVBlgEpHWOspbMCN8p79Rt0PRCKvoXeouV56u1TdD9DsPEol0P9+M+YHaPsF
hfABrJCgt55GONAi/qSeeVEr0lknGeryPlLtWKj9W/qW7kMGh87BmGe7GMPyF/VnaScNDNGv/7ja
5i0ZRCsejMS63peJ94xDSSJS884YGnoduPADBmDpgPgFoNH38+xiJZymfqm4u3o4IySe5+xwB8Xr
W6fs4mYCoElopgIgqhWS30r3gk5csylLxZJCA1Nx8vxAgiz7wQ0l5DvVcSTbmWK8jfHxqlAWl83N
NB7FaoFvsdsStBoi/xD9FI7qNHz5pGbWSfA6zzSrn4KkFfJuxy7FOGyFzg81XEiyLUiF/11r/JIU
abdfGnlBxyyp8DXCrx/DhThDUYwmiNqpc1uoNQLTdEnXs7jCe2OnergVUZtsmUIh3JVvWZHSISSP
kSw48wrVPTSkU5kLXSkJYQCgMmGSypKxDkLboAXLFO7X0hadhItbVcjf9GTwHJE89BpG1k/GKg+L
TstbJfyppSQw84NKSBV01XSObfzqo+e9QCJXcmPjvU2VP0sOy9SYJbCwVyKH7Zhv1dGxUL+uN7uE
63J+uSiO/3c8a3qAFpSySEERtJ9TvORF17KR73I8/s+2MA3cxhOab0Lk7fCXR/IK6etaFOoiQHcc
PE82BrAT9gkMRHYsPJZe1tY8eFP+PkdrmKC/yhDvNa0/gewF7vCD5CRDn+F1VRhq4T6uZeNThBqp
RD6t8z1JmMUxaJSDpi/aRPRgw4qUHQqfN/naux6NtO9M19233ziC123L1t8Pe5tCFsa2I8gLxrNG
hoypwuj5pmtL4Cw69myu/3TB7ZSNZMvhK3oUC/mP7FverP8Qk3hzBOFvhKjjO9bwZFmQEKvb1RQD
vgj0gAaCgbTLgbcVSY480h8i8ru9WOFzve1YECduXKdOdgJxWBmODyLNTJupwbx9cAxfgkYKfK92
iGpzliDmX+kjPEU2EJEKd7v4Ch6Zcowg7Ca9lEmvKHhVZY1B6qw9f23+OP4mE9T2Ukjgzs2r7lwr
ek6ltHtcqP7byGNvoWhAk3HJFMaOZDPNzfDeMbZBz1BHQmtwX9Mq0qXy0rh34yEqbVimmqgSXLtH
WPaMGq7sgd25BVXOFixGvZyG7be7hJhesnj1r0w5Otg3h2z5Mgy2ccQ2CVLlJSl7icdRCwgPGRm2
d6kpYWroVt9w7KFiTLStOHuHvJ/c64MSkfYffGC7ROqgw4SxBctGCm9+lEQtX2daBPvqb/OATm0q
HqNdb6AvtW0R3q2JfgYU9fEJAMqQmduOzEmRSoVZw4OiIXMOFgeAUWUz1e83ogO7ZHp4EikMR/5q
16BubPn8bvhkPvMvbfFbrGV/5AzXDr8HwM/CZOvU/73jEvPDWyo2CfX3nvink3XX9c/c089FMQqr
hNzKCF1RVV7d1qGmuQHlgH5a4+QNhcD8Wx3gyAjGpkpIomxqPrizctRXxoeAPMUClhpTXhYA3TNm
YkvOQWzvDryUTyoQ4t864xXrPp8r0YOqB5t+b+clmKSwaA1Eaz54fJxVjEehEQJSeYf1XhjA4PE4
D7jhLVS6PHrC3qbIxEDQrBEI5w6x8YAasAMNrKdozBZs98oakQbF2ri08meABOj5mpO8emmMvGT2
654d02kkyZaxq135k2KTFbEStxVmknRvQrggQAkBuPT4ocLTSmf6kqly4YS17Ljr7sFEqgm8Vhdb
3i2yvVW3kfXlH2H7Tq+f0PUkKpXIO6fRLAhy29j8KF8lsrGXqqkgSknkC68sSFSiMXEpBdtLx4Mg
6PQkSjysh/tUN8Euj9Q3bR1oYBKvxbIa9KVQiAdgwlNjCm9YGxJMwqRMdcEbcaxqUiVF0u0o9kC5
KgytDyKdoEpR3yfsS+AEzaWxCFa/TmKZ3cDzqfAjGmcGZGhTQj+r/nZ2RSWDTH92pixSoHYd1aHo
kI/aj77xwAwBguQh7nfP3Y4v4vhqFqltoK2KI3o3SbezOrSUU7G5vZQhYjufgQZ6oE6q1MVl5rXF
u1NgxvPiPvSzwei3UdGHDfAvnrZOs/VukbetY4HfLqJzf2PI1DtY82MxGUlKUKUAqolakCnlJHQL
9zfDLK58ddDIxHBgDv6Ak1VVHmQN+e9LCpPzYIIwCG2K3/inHE7f/2t9li6hjB7nh1ymGwtHQe9N
ldMuLuH9y7x94DytiJ2B+fzoJ7+S0vb6GNwY8L7PfYZXfDrroRjOFah25MP3qydzV0ivjtM6IRMN
5A4Q/3BXKB7rGePvmK5nES/3YrvWGrNYXbvX3KUrFhSqWmmIP7IwsIdWpi3DNkIRxRletD0RJY5u
ZPEQHB5ySvR7fRqes5hbFEYwivTyRYpmcBKFPSfyjF7cOwlpA2H9NNUUhNy3IgVEBU+REbwzeLz0
DuhLTd1mDYREXJu2VT169tDZHqINAx1nyK1AXpZ0b58sDy0TSKvLQS27dPywfehcvxfCK12E4zGX
lsx0GRq1se8ubBWOfRT9VpX3QDz1dYv8xrbPT/7n0dheT6GG/oPC5AL4IxC0SG4AarmqcZ0qqCvs
JodLH36JRYPycxXzu7eHVmAVoJF9BMVABKu5/rdd3JfSHUD7RZy6ctyRRst0sftN55HX2XS7sTH3
z5KFIqGUmW4nRtakEpKa7nLL9szJiiw3Ipj4L2sv6i9Xyt1ZDbVkEI/AqkZwq9wuJDsCfeEPKZjR
CruMD3qeUvpULUpt/AV9+BEkhIUtI1nJMjxB6TfX9AdG5Vy79FyK3Qh3eULFGmHfVA5TCs+ohUkH
JrCzNUfA68mYUdyDL5Ddtlw/arVVsHzXGMo3bQmizQoAKfhhLOJOkQ/AmOGYFjmZlx0qVezqEPCk
54xcJaMb3w8VsqFHvnebS7goVllIoXRBfMTxuOKOKlPfgmCssSxlaXR1LSSQIwlr8RzlyKbWC/sc
RxWywKz87eWQNPl1rF0HgyqRr0BQs840GWju/cNuqYP56NBZs8FGUHjBc4sxpB0DgyFmXn+ZQQrZ
3DNM1P3sY0iH5PtH3U037cye170YPm1U6HKZUKtKAkcn9igz2ANDC/FEZ4lWQNGGOf2Bx14d2iAi
O/SOF6ZOkP6+COj6RPn91vbJevsRi3BxsYvl9gPsOTa0Hy+VShdioO3RAhZJM8lhNsoiMleuhHTv
gY9pPle2Uk7NljXAb+H/kbX2qThxQhnXF0p/Nm+/Mc6PUX2fTUPBdcVEoLVD/SucqcntH8/KaXDF
mIPvefNkzyLN7fNFlk5B0p/hj+3/Bcs/CzauYu/wijzUrhTeBIQ14NyAQ7YjNrS5by7xCNcfjyGf
btG2LceoOrW2RQmzM9r0RB9r1QGU3l6zuJxGT5xNUueVoI9natREI8HLxZmv0ci0bLYbx8NZAjHQ
FRma3W6B6hNY77675J1HaAF2E8Gc/pk3dWmUYwuLCqbcDVgFRjYezvAB/rKbnQZNMv+giZlksT7a
3ymM7u7RUqreVDjbxBT4ofu9Skojuj/Z4fXrebEmgCi/vaeE6PORiadTVF4mqyWJyHolujjtK4KO
+AJx3trqdHxmX97buFmG3PocWQE+vrabtWkPhZnvVcWdhXfUbrp7SuOjPrZ2A9fNKETzV4VpJRGw
zI3qLDwePy4gFskmA/gvmSSpJzbnBZIZH0TbH6/XorXCqAhAIMZ0uHCAPoNWzZRfmDqjrnDXw/EU
/I2w2neBoRIbE41z6S/mWoi2tqc0alSajeTqf8lOyCG9tfWs5x4u1h6qADnQkbWRKvGPHCh3xCpu
8p4NFWDps5XguQwTQynKO+pQpVhrtET2zv80uivvI2F9ZsWQa4takbML0/TAYjBAQbnpTitlnvXT
aCQWvPv7rggPmf5zxUYWEQX1aKCO1zM5LlkQ5D2diaTjQBakDx2cNrveHNNrlgvPsWnt8HifmZ8s
CTcMYVFQuSOWDg0iqadNcbTcYi6ASKWmcqfogDzCTuJLepijlCzwOcVJmQfRuglpmViKtksDCC0x
IxMgxN8UJ/mq0IUK4xf5iFxcQRiPhQWu/Vfox7Wq0gGTA2a5YYHtjTO3y3WeDaORiXJjv3OI+w3u
YKLMQ0gfv0af/vTizshtTySy0KoKIKwIgE6IsXSfHSCx0/g9Y8CZG1BRJQp1zWxTydu2knYWlnHX
qeQSoDortDS5z6SRGos4HcqWSWuMKj+X5x4n/IKDB0fKBQ5UpC1yH5nhYSFjMhEXS924HWB4BzfI
HqiflGRmgrx6gsMRCxoTgvNDdfhzViT9qF81JtTti1Wy6/7FYzbGtD9+xjfPend18qX3zWUihggE
1WEvGy9y89KOygoiKL4Pq5HU0L0oGhcE1WV/1woXojFnG0guld0YxUnbaesaEuT4u5GtqWrQvYFX
6DNG5YMP2s6a48yHRStYdvEOYpiM/yuptYVeFBBfsGs7fgz2wybuzPPBo341tK7E2WDiDWaaomf3
KbiSftJUq3tSFrDOPWx+QG2CDXtN3v11Dbza8wcdm8O2og1Oyy6zGhbT3gPLF6PFwkuphCM9ZAmp
P6qgVAuJJAZN/bUDqZ8UpwwrwqAzW37MjQ3FqYNxxDqyFcS7COasMnsiVWDegsFEDIWmVZFAnTgF
aVhkGU/71UIumxETm3CfJ20QuHrtgV4ZbewTrAoYmsUgSqZw6GGjR24hqgIZNFXZfNfSMJfzQMAT
bT6EicQC2L4dVQyrGwDGlzL9h3MdUxSVu/7ODc2jzcyR3+UND0wprrN4ELfwMBoyPwBs6Zz4iuK1
IRQtDtDHmNmePfZ9UM0/SnoWD1r3GezzKicDjeTBH5UgOSiWn0jJBunqoN3kEHLxhyjnZg9CWeMa
xhM9w/Q8zOYSosLv/W59aWRhvkEWDsSsHH4Joh17tSGyulezcVYeFpIdAonosy1U+eCq4FDvUHKb
tzMnippa7enpPcyiU6R+VPMIFyewVVThRrXztCU5kQlAydK/enT/lBoGQ7JwFjtOjwefoGY8dqld
wCtNBZkrMuot7AFW1cLzBME9kBI7OdE1CuB9zJhzBhTmUqUsT/lSPa0l54G37dOOZ6GnfOXKyEFb
jCgwJPrnF9TxNFeCrBf0SyC7S35h1n6xTcdkexcGAFT4E9p1n3Gz9rciyDws7uQaboU+JCOsUO+N
iSXJjzXAqBUsiZWaCSVQJkAsiJOBwQpCjbIRkzWIJNWBN8UOpEglxmssaKVfQYh9jkjU+GEDCuVk
4vZnWrrsBcejC3thG4G1sk4YmwcEkv2bVMe8jNGUy3cE0L+60cgx05fqG0JDfRXoooT951Rpto9G
rRTc5UO9MFCukRC6Piu1Nu9HjsHxCrlUmprw473W7k29tIBW2m7Ljog511k8ea40tKjMqh5Atll/
1EymYJNH4yy949kSIfi/QguZ/OORWWp/H/e0AMEvtpxsc+XFSjmVmlgqa0G/2bE8NtODOUXX5ZnZ
cpSHEPHoroFblM74y3E2Jt52NdhRMEXYs0W+SkIbzDHXxK1t+r0owZVjsakOQpHUjzgdHoTG2Aey
8r5a601MyXmVBzxrbEWcJo6s7NHlhCjxu5JJr2SiAMgzGDHrN4CpclmcTzG3Ty+ByBm68qY7Thbb
Lq5Wc6avTlpUq/Q4zbUOr7NEp405WLsmXPna8Yk/wX3//XHx+aOth0ImbUuVCnfd2XkrYo/JF0Xr
M0Bao7JbFMuDJ37H+cRj1sLhvkPieMHI4oOGNUPQG0GygP5wduuyEW8Zh1HkUNtl5B5YP1Qfs5qB
KA/aNE+XnSgN0ipi3Fz834LVGO8pRetV315gVUkJuAZUVveCCfAxxrOmHR6X6X4hP64tbB8mpUH0
XkKX1bPSPiylE81q9++o+5dVI/BmM9Sdb14bqBqqylr26wlvKThjT7r5hwNG3Wdd9oS9l+u+Nnbj
45MT4RFOOfD9vMeZAKef8segQiQ4hq9GnYUKQtZUw95yidLJJu7nU3agZ1Ygxnx11j/NA5cUjFjL
2TXKAxVBImFCyR2cDkMTVwl25kIszC9L7gGShLoSGJnwXSMVLyucB3vbZxOnpLAbQefUV4BMjK8S
XOeWC/lcQ/1kTLDXreiKNDdlxuj6cq48ZiW6vntCP7YeYgE1riOb5kHAuelFQ8JtOOgI1DWxudsq
9cryoZTP4SV5WvRk9VHwh8bdpKscnwfGBgH7RppZB9nCIcNofaCGSirrfj0HlOMrRzEaciQfPjj5
I/iSlnpXxbi9jZTytAEZrdEKc2qYXL1PzXoe/F9TvqC0qwB6hiHhMQv/f0cUwfz2O4fee1yO2ygV
sGyWaPOYwVuO9Y60p3V83Bsq0w5d8En5BSLA+J80qAkebob3SAmYg9gqpntTpbH4qJW0CgR9Barl
L6/36h6Dhlud4wu6t2JDz3x2J5oYvvXOY5za4L4YbaoRnayDhYBe0Y8ItCE0qgSoPQs4Hjkq+l1p
7ekZwX2mpo1mLeCBFlg4okjJdXOBwPQAL3niDbZZcVUQc3rthWn03p9AM7g0RLtQQqBFfcJSpbTt
2vJY43fBAG38s7I8erKgBS1mbVBDu7ZYI6eN9bcB/lS4GPSL2a9RcPzmkI9xrBC9dxrmRREcmi5x
drXekGeGkbuZvXwR24G3wwOMzAIytfxOaCIDna19uOPdbZQe/TBG+/w5vUkyhqLUd7qOqIB1j0Iv
NPW7pfzuqrA00FPQltu0+OihNqcO0w+/WQpAf+WSujOhUjaeuRJNo4kx9m3oQLo2ReuP4Jx1yCcH
S6JFMlOY96LXAYOFSd4XJfQXHFDIbL0GevKD24N7b1C/9+Ah6jGpFTY7NXuR8bqib2OjZdHeDLE4
/oZWO+ADsfFpTbcezvk1qy3puqNG6Ytm8W2x345MqpNJULQN4wnsnKzQCYAMKfbrZz5ZQcRVwki6
nDz7pz+/ORpOpRqjYLnjLS3a9fhnXG3VLR8U0gi2WN7LGaBYbyG6BcM0D9Xj2r34xBa9Cn4/Iv4O
mWqdDamAcCog3YtPPTlkqCd6oATfFCtbEs592dfFK/dQxKzHIVvmzSxAKZoi9/FKLCYyJz4dXZQb
KROD+w6/61XJmge0LtYlxeldebCjMZia00x4HeRJq0yfY3+rCHsEP2veLYKKOwvkg2HA0PP2J+K+
6QPGXoZq1tNlQIXS8VuFBoaUGnRF6EqfPIPty3CHsfuL2qL8buBhP+Lv7WRC7CSA8ncPAbj7E4g4
4ORnp2XSe7GK/f+T7ydn8YUuoJO7SWwSAkQLmwuTV/XENWmXgQaqYvtUDgZwLebdSeOu7v+6ormy
XFR81FjxOYRlqK1NO/8Zekw1vVk9NqUXhJcNaZ1CBBJyNdEfZRSWB3xx1hdn6bURjvjgFRUymjEw
AiJwptp2Pnpxp25G5HJXXKj80ADcW1iNMJPRbxE030WSEBa07xdW2C3N84WFSAOoGQ+df/EtaMuZ
JyloqajReTVlOqE7IsZ9GrrbN2ZlvQA/iOB591fSPc+37fHnP9ThHJqi9rEOoXXgvK7AOs+7gi52
4i7H+PKTNpYNKPIcJmLRhJlTN2OSANk3GZTBZrBJCWvjZ7xR9nZcbAgJL3O2hGhFm5/90Jk42cIt
UrQpknv6owkuH4PMOsKCxKz627lrlg59rktS2OZIU3IOIVatlBLNx/R47jx/etJ4qxDsJkpVjTXt
ntbWxalAaY19ZGHUlUr1FJ9JZW86dvW+hOsDgVBm8zvIPQ+vSIxthuzF6zr5IgjQL9LYh73yyzlB
z/u9+VD5nFWKdoD77b3zcc4UN2P8EGzHH9lCYHab1AE56/tiph13oiUg84v3pWr7utAsM4ZrSPKg
lNqNiTzmuCzlKxWcBm/w4Y9gBo3z6LyjFOlkqH3COxQPAjpQXk2cfY10JBZhu4Vvep7w8akxm1DD
KM2zO+rbWzRN3iHsK4fsu/5P2H85mzcXG5v3Fv4txpnBKBipTPm3fq8ffBvEmEJ5Ciua962dqWgX
vMoSKKPARchT+lFL1cL6ewpTfU+hd463CeVkuzDjsQYHxSnVnQuh9yOb/cvBBi6Vv/tlj0v4d5Em
qfr8v4oXBZML39aqgWGg8Znwxi8dKPfKNaGrH+DrzcgO0Dwr2J+4PlB6sFWaR4gTl1Rlo4dA0EqN
HW2k6QqFYI/iQJ9Hv++Ogrl1SOMhCQ/N0IV78QuOfMZDNZtAdGMur5iRh2b5tpnvSMOHhfu7gOds
nCwnjrsjZuvYnchSBgAOaGeQwtwz+4mKjhYVoQ0UTJg3c419NGVUoujoEzwLQ93LtQYM/aHiFOzh
XKJ373QSZ9deNYIJ7gwkpGkQzdCRCsGI/NCjss2VNNq4CNiKcojpj9RjYNPgrNLu89bTsfwN9w7G
Hmqb6jaF/N4T1yNNoPQYAM5cBRk6xDCscw5mMgTfZhC6V2jHLGkZ7xnF7/FeuGNIBes3I9B2rYBC
1NcBJis46MtGdkgr3Cef/8mrx+kTTRKzYIXokwprSEFXb02HgO2fjK1GCRMHhHgbQcAeuF0eCq7H
dmWllI5L9aHiYnAZS81pPT87Jlze5pLw2ZjPeVlKZSqssS2tO3ODscCG7+6HHJIyWiRsbIioM/a3
crRSzzRSKOpe26Ir+9sgiFgko+VD4IKjtLBvqOBvPIG/ZUCnvGGADsG5RkrxOP/IYGtgM3wG/S/V
YpSGSBfAku+3kHwjoAo/O00SGp7WB9LaJl54cmtcxwRNNinCAK+803h4Yj7BUvHw7WYzELeZAMro
dM2G8/0A7xbG6RMmEkd+qOYlHdPXpn+tkvF2WeKR2I7IolilGZ9ugiuNFFA4UB3NJcybYicO8/xo
bjbrdo6Kj3hbNuW2Tqm2SfS7wc6lD2gCLqFw0g/TYW/UsBwcwo0oVtR4VIue0f8VWr5AzBppa2rt
MHh1DnNJYcDDpHK6GjhMid93b8U94SoCzJ0CiKwgIOH1C1DFAnrlEIcv0NldvW1YvgCewi5/8DBT
HeK5T2QPUXbnE5dlrMau94/TgIXMFYW2j741dKjeKIwE9dihYbRc6Vod3O+FnIWyIHs4rr+cs+8M
195RRFB5R+/0wi6zDQQlzh2Ut2iMJVPmbca80bz7VGmoiZAk/pL5vpBabm4g5s6IObprlddNOvat
0nPMO0kXNR84DlWgMbPcAAlprNrx1O7M1fd7Ar9bKcWCXjlUR8SJ24u3Q8IqO+PophH58rNXLUfW
pF7Otd80cBnDU9/Hv8bgwh70owsiXUnLQVSwYZP3IXihcrQT71p98Jv7Bl6QNjxwsj8Ne17SpcMD
sDjO7bchle/F9Iq7m03KGoLnaHeqqj63nalTz/XFPA+ZJDEBDHUdLC369czQ3yI3I5gMGEqyQeU3
CxC2FAjRM7H+92/T5dmiIC+A5aOJi1glrFF8Z5jN75E+dMJN3E2OZlN2MwSnk1QtgOrPpOCWbY1d
t8ta93C0/wBnINh13yJQpQEyTqPOptsAs2V/VOHso3xGKpWt3JvuIFB9Q5oEwR60gL6bARfTpfUv
xuJRJuyUs0XmeAsca/KmNOvdAp/iTCdJLZl5ePoqU3bP9d38L7pCSkGUhHIqrSLGnc66sMYjCcFw
1nYO89liqxeLv0S9cr1zX9T6QEhf4mc8Qd2X1BV2RkQFvcfWYU5dxcY1548XpHrSbEtuoXmlrrU0
OxTC/sBWUebJvDwBD232zQQ0EolcG2pMaTCoPwjNpoCaMOnqyfP5hndTSCaxSyqS0Zckbt1RPL54
gj5WbVg3q2fy9h1GCxZcXdP3YJtOqv2y0193m1y1d41sdGBOnkOPF7gA59sRRDZT1RZgbt4RF032
Q2JAlwaBw0kuDfzJPHp+A3Yn/91IKpdE0HbPbk3YO+bEMYCYEKLJIJ5kHVfgIBx01PkYmdzuIlfs
kd23Ey2GjG7TAmY26e2vV08oQp4vkuN153/odjR8qmSPEyqgsmK5TvUoCGUfXNuS86O+A6wZp/RW
lXZanCMrXGxNj+buO5yFvDeRco8RnQI5mEXXq0twjAtM6+n2+KV6TrOqOcem5bpXO6PBMZuYbmga
eoAgqeF8O5qgRyzAx44ldXkZFiwwhLvUnxRrAHKldYVfVy0+0i3k876R4gWPIPm6/BKwil1Eca1R
5P5rEh7f5eScaiayV2Fb6OAHKO3WSAVqnYEs24DJquobhNKDIO9FRmfSME17ne63V+crINlqGB7R
27beIpTK8efG5lAve9Iy/H9vyepFMvGCQs9DapDiuR0V/RUMD26I72Cz8OCXYuyPYgeTigD7LijB
A7spRdQmbz2ioUSSokXeSa7watISpJDKukwRpCmhJqPz9W5Y+6MSux+fafFbT0mY040O8VuouMJs
ivY+8ZTNW8Ieb9D9QcI9EwdUoGAqZE/6Ry4caV4SWjXO7vvnwX0ogcoNXQcrfqlgIQ/FSgvbzhUT
1M9bRD73N2+i4KkCu+ANwpd5lSLVCdE5Kwsg4lWxZKAzWStzOI82+oThImVubfElJNFqJ0iDZCrR
07WhdZe5cEkaVQszp/qiPxutk/s32DDbLPWQLRdztOpREFUjY2S+5UvGWIoIYywyiEEVRiITUX2D
cgzE2eNEfR7KwtHRnPA/Edq2lUQX1JAeH9dn5wg767Wgy0T07Q3+dtf41qxdwmKwefP3eJKP7RH9
r/0cHdVdmEdqhdO/a05RcaeX01MtqsCcN7kxDK0JlhxFQViSd7npGNYMwlxm5tuof1c+KR1E3xHk
NtRczKrEc71nL+pct9ftH/UcKlH++udFFK8QPoovIrx8UTKS4Usr7IVggG6kvYOE08nrtim9/y0f
EzzNCODMdoYW5I+WN2ve5wCvEylnh0xD1XQ1hQq7BWJAmWv89/3JsZw6V4h6dUxXJehXBodp/fE/
WEBjctU9HNFgiYHyQufXqYpWe3Y/KuEUL8o31j5Otib41hS1TYsxqrJTt/q71pGxrO22BhoQpTK+
fABkC1mP2Fh5gi7OJeD0K1Tcf8xn4FBxkbaNzQ+kwn7o6YSZhCl/X3trd+2UIKEVK2QxESjXE/8D
a+wHBGcO9rlkQ9TjBkEROaMTncSnsC5BzpzTUG/cFYabE0quydJYBnW95cd6WfkxXmcjd3y6D2m4
W7aa2Dtl7ynIIhNXUaS/aK5qGZbFLIb/3k8LscPTPT9qbSDVnAzZ/tweqQ+VbxsCBmVQAVFMW49w
+nqRFmj9Vz/y4GxszGH/KrBtZrzhTu6OcPiEG/nrLeRAavQkx9YGwevadoGYzHtclvlOEaHhEg+s
KW+e+15v2HBRPoz8q1R7uvMZn4QXqlFCKtI3jDHjlL70XBiSdQKRurKhGsJVioXRuPPeV4azpbjH
SMI6kwktKkHibyxQwu7uD7HC9o8vBt8I2fc2uGX9rLtfb0X2njeAV32BdAEPAs6ojaMBFn6gHuju
cztFhI3ADcmCJZefpIVsZ2a9jRwrV2g5nk814QTR32X6V7AS//GP7sGc7tkTO3euIWqn2f0b4Vor
qm9xe03BrenA6A0xMhhA5y1SMWEp8Xji8yhxjyfu5KhE5dk8OGb9jBI/WDn/lFKUf3IRZvBlgjDr
B3EEPbkF/kPj+y+wO7feLbQ8ckZk5jDVRvsJbpGOWc2lsRZjtbvWJX2SnpohN/iM+OK0SQcuy3+N
RTNY/W+YbFsCjVWTq5XEnEWktVy9RKrw8PL3qdvZR8fxQlJaJs1aRZtFgNWOXND5/iLWowz/mwYv
xcKAW+1Q7Dw3ZSdTFpTKjTthLq5YtR4M3jgNFh0FEEz/hinfjOp1WJfaysm9qLwRyFdLlWGATiLW
AOZqDnSkkUk+KY3+vUDZIlw5kU3nTggLjeYs6w+744iTj9zrQANGg1oX7MOuaKU4pKO1Mas0ALnG
fM8pwj81/XnzXa47mRz8CIh3nZneqr5j+PviXSi0cVXCzqd5DS6PynTgV5XP0yzispxHF2+jSLc9
uBCQTq/15tQbnKTdA/1erb/Mv2MCUH1knCui80zB9lNkReZdealhEN+vU0Yjo7kaOW084sF7grty
nRS2t5dhEb4q2wtvrvVTLLrDEtjNoDMYeSNQXy/CpQgtnYeW3bf0DOH3O9AZ/TYHRVrA4OxXp9ap
AwuAr8SftID1CerwErHgMqsMHgbnzDFrBOWuSgFX/Z2VsRjwQ6yAG4wCVD74f4VHAW93VHH1fzq7
Y80m2qzemFTBHGeLqDMlUup9vT4zWtMFQMEH1X0X+YLQJOTABmHBbQ/VAvBSUsnUh8ju3Uhn6uLn
iM84TZkCfKasnd1BHoAwtjzUaWf25mutHxCgJ0+kGzA5E3ulh/BPU2LRDj8zmkqgEq06mNcgD1MM
XXjO3bSYTNCsSOfoINaLd8cmg8EoKJWnJrg8zw7reDh7p8jamTvW/bANQEPsDmQhNflk8+SIRugD
JwNgAsF3q8TXdiXRFx2mr0ao4NOpC5HQc5yJuvEWl6uQCttSl0fJk6uOjmtnBqnJVp5lcCGs7QrZ
y6a2QrV9BIwAAQRVzZUrQ7uTdwu/utisdZJhYujjjeQlEuJotQcZAZpwxBS0cMhG9CJxSvICARWy
lM7fhz9ycu1zp6bqmHfq5vGbmJqw89K8MwKbMWJuevL5hMJDbMdOfM2C2N751DV1FK6EZoUX41e9
y/LroGbBsPo8kqiqLH98pBfSz6dFB5lvKS5CEKAOia/K+6PvfGtnd4Ex13HidMADUNLiAUmprVRF
3LDSWEZNqPUiyLkEoBHXREdE2yAi6DuAVjX/GGC9BrwFtSSWCWjp7S0DzGFzxIaGJSbDt/8n1TpX
Q23lxc97jU2K0fQBMlYDUMrlcKxcyrCviNHyChbVuwGXyNO6WGkukbfwFPR5HF8d8qKgktmcq1lQ
KTHuo0ecruhp4DYJPOpy8UEhEZqqE/jkzrR1NH3RJOvNln+r/Yb176a5RTWMT0xihH4324YDxiEK
utdr0K1o1sXDXpzEHiwL/+/W5If9TpyqKgKY+gJsZtdSCahoqTw/tLM2LpMCg8d2a579z9Kwxeg6
fCNdCfC40z7ExSCkJS4ErwNaPhBOcaigC1B1fCwDx2IRsDdRRj+Xj+fQiyuZr4F2WzSXjAQXmMGn
hK5KkXPKEwZHbfUvIBqeve41DSXXIfYHORknEIPCnjIBnPLcb27iogFVsGKYiJYNaJ6z0bwXMROo
5mTfNy5giOLuxj6FMngL1QCWN5WV5UtKRpXWYPagbJ4rKyBoznoQJw1ajBd19HEKUpYmNMkWKTms
lcdyY8Ug7IwKddRekFUyBgjAbOrI/IY6+8yA4ytodYJz9O0UhkvOquG+2xmymqaP/LJ6X6xPBBv7
I16fLDFVMavrwA4BzRvT8gI5EJ6Ufg6GYypbx3KCTJDf229S0i2ED6GCN4ZvIpYGbdEyQbppuD4d
A+tcPWURRCrLHUnOwd24lwv4Qgmp8XS3hKaljcWPpn1klAs65h7DO9JUghteTndEmIKcfNMEotZb
ZvwwaG13L/qvhi1KbFFg+EhutnX/vMWOnU4/PjO5Leroc1CgOQIGBMiJXmOqVvrh0mgAHnF7iRW7
1j35C+Mlq1KEJYH4+9tpPw7BjTAe1jHzwA0ULDkKfypOVmrCc/kyIH0/5+k0Y9uPFDlH+pTR4/5G
hrk0bn92jmqTAI7F3gB0j5yYb2vSgVCY8XAM22PeCVBt/ioQMCP8la7X8JTVBzHK00Ce7Kpps8mN
XLWqwWMDU5o+gjqbEpIFFmrH/bub+z4rPFgat/i1lrqxYpJC5SY2wJajcSqfT1cQd2Rr+hDjQqpR
N0jd/48sAL5B54aFrO1QaySCVf7DsGDKVvyEeNq6GEdJ1YWZW0NH1BvaguBJJJolrvPF6E42fX/m
Tacw3/g6h8dl18zSkX5FA9AYM2y6WahC/b2EyuTgcpg6t5aPQdlsXbE1t/UN7ruYmoIIBnsKFN/d
K7NzXvJZ5e3HlSM9RkQshNvL5W0R2vVom3tw7CTWbMaWAnXkdHHwh+pDJdn9usN+SPNMAYG5Veda
e0o7Ylz8/la0SRFeumd58PrvzsM2CjO4JjXwAlWhP3Se3L+SUkzgHoAbXN7ONXOptQajDWkE4lf1
MrbsaBaCL3DykPfhjvcGBhAvTiFHlO4bUCcqneR7ex3qQWmr/9XIG2yv7AP6rZZUb71u68OJC2Gk
BVTiI1Tfk2jnINfwgCVUKGuZE4JvdWCQkmsWPiIS2jy2/GDhdBdl4Y4yYAB5oA6TVz1LRSD7kTMo
UaKkZe42QxwcItCw7RHvalgpx70zgc2Omx8zsSrWik0S8nGSq+MG3wGHPzpPDfv+vsc0NB4XUnhM
JkF5a5rdKNv+4s52P+5rhYNv0WI3s6Wj8wcPn7DiyaP84JVM9si6ZoA0c2mE3rwqcA1rOHQZd6Hz
BzLlfUOe7zXzSWgRzkJA/AD1cXzxGB2Q6KY4qMmu2HTVo0H7JN88coc5iJab7IYpzkAtCuCRNUSK
BEirL3imaW/yPy6af1M+TzKEB6qk/RK2McGDW1j1NDY8xDpjqP9FrdtfkgEVvRAzIWEAU6yJnvXl
o5n7ExVVO3fFztYc063zWnLGFOx4Wmbwxnx3xYhINMukzQ1clAP94bTwbjfKhlgOJdPlhllTim6o
JYBfTChPqMEMGZUjRawe/KMa5dubxBz09qBGqs5bvayFuIjXyL2WZ5G/xuADQ7KmCHEXGphdo3+i
qMxGTo7f+4wJEeafyFZT/kHKcf+yIoDOD5QcbsmjJPIeMqTXZq21worRJGWNytBOrgzOtH5wXgOy
4PPJTLHNz0m/hrWETPfWdyuA0rfRcRPjlwl6K+mxwFd0X/hHdOVWtxIA6Q1e8WsBP+qII6vs8RQQ
5bvkEvoutOkLos/G3sBrgBfbpht7NrRiEsoas60d/As3i45uGoo6VKZ4B7dxNHJpKwOBwJ49RDOg
+kBcXoN7+dNTw6OTVvBSF93JYBs2iL3GlJ7gfKITfTO2xo12YUPBQSd38xxWCbJdXrQtry/BnAJ7
9Y26hBbPPvJroX5g0MbJ0NhCxPEvasHZKrvynMduMoH0MUYA61j/SAQFQXEGodl/MerQncmPFUFM
OhkQV6195NPHJN+JQ7HK/1xO/nbrS5m2zA5JTi0OzrcRxcQ6JZDCcrNJN+hDnQkogN9dk2g4hSrc
tygGlRror1KhW+6uf78BheF0ljQZzfxZGMad6np0I3Xj5DoIZvS2Y5dDWWo4rEuPhc/Sd6G/dIz/
cN2sv291Tb2p2zS4sZEgbXWq/3AX683tTyOUGdz8YNE5eziAGTJf7epoUO9kXolSz7aDjEFdSfb6
A1o6nNDLkQgNqpxKVC41oEb/55GkxIkabwd9DZIg2aQQxiJoaT1fKwjyUrX83isCdBcoepX0MqdD
MVwOe3MjRyDts5+bpkq00eRXmNyU3Ly/1Gwg9ywRSIuv3k1aPg7kXV1Ublb1PD/FtNBSF9nxfygf
kQb8MWft+kOBxMr+uYtkadBl5boSuBFhqDapYOoPdyxsma1BH0DtrGdZgDKQdbr3iZQpZYy9+1UQ
wR9JBasartZlYIbrhiCwf+bXpTd67vybvt7YahwBZNmMXQrngWacHj/pYN4mw8W8dGVy1r+rrz9h
4FTLLoa93DG0cz7HrfsN3v0kG58G/VD4GtYKIjQ71uYbMcYfxvq0/hWmHlf8NYoP2IgL2VsvPHAn
H8m+LalQawES36pMn5e8P521ONLbYlijMpCbP0N85ieVkQ4ZeyPrcbt+aP32RgqrJLCh30uos/9U
4CEq7e8WXSjasfP2M/uVq2bJ/LZi/nHibgreU9iPFgwGIy7/h908JHUOUJ3i6Jd3v24T6+s+qU5a
b5AU0v5tMmD8aMFuFNoZshLqABb0JmGGxDez0Y1FlkrpBf3j2Ikj/SZCRNvATmTAtFY7b1hv4YvE
k+unwN3K5SofZNbebqC1LccPdiTO5LZkSwe3/MFKOomZrPoxppl+0YU5OOGq5aSiZEdQ51CSYUsJ
kQFwzBDRzvupZ+LE+X1cJFrifkWdkADSv8qRJit2dDHrA+LOPWSP/p75Vn+yL6dLbdNR9ra+Bw6s
kBnZ+46SdTWR+nF8ab9FgVkSzPWHJlQdsT9FS6XLb73ymSQg1CM4FOcyczDnNYKsr1WhC4YGzRIe
fP86fC1wUsJP5ZbLjMaCMS0xRG7alleAA6jHX7KfnUSUs3jXcNdkvKmxdzp2VxmtP5jsoZS9N+2/
DW6ZQNquRT6XHzI3nOEcrFSfzQLP/8oPgyPIWQsXxFoqpFH7Pnof793TFxU5Xd58vfA65zvqU0o5
5HSW7wI8Pss0ku2dmU/SNxHAqutpiQ1lgZJq5t2HJw+dXEs0SLwZ5qIiGtzSF1ApCsaFS7B95VGt
EVCpI4nujwNPlUsl7avtgs0OX5TD8zai8I8jqFdjcrGrv4GVHlnYBEWwIdX0fZ6YR1v4Xr3yL895
cVPmzfzO99nFEnOsLZ2jZIH2IOXsLY3NzTPOxq/fJ0XwxyENKRC9nWImvYmFXxslE8a1EHaKdK+u
oWaWaT5wRlTSnqQ4XG0UZ5PNI/tKsnnzgA4T1Acu5BkJzkpsBuY8+62dRt4wkFLMy2FwTfuRXCbz
hGTUHJogIJ2V2jTz4SiPXNIkPl0OKaVzf4zf4BUN05kkbRbYI98JhmZb1wuVWpTSvD9N4TMIb3XR
UNnihW+az12eSkD38cPl4mVFdi8iWWB1Uld+k5VsEnPtzxba8uSijPuwpalayMlRbbY7EkDCPm/2
riuqJZ2LIvE0uEPICZDWJjjzzeD4tkON/llghqTncRElKTq2o/ddyRio8zV7ld12t3//bslIpPYR
XFFpVixDKKJ+sqTpV3AwND3QJUAnU1f/MM4ng7fmx9ficNGBs1TJeNaq5tGdNgBi0cR5jK4rGDLe
Lz5nXghjidoPsAmNZWhrq0v5YjORGrv7VT2GNm0y1qBCwcs5e733weQ6F367DxYed1e5YC2g68z7
x9iChHgcsLxyZpiMqRd5yMGd/N9h0/aEi+BycSX8R6HvAVkFUeIu9cqjYtTaIlVBjZQiU97JE15c
ATxUlcdQKmiqTj1M942hyVafTpPy/8BQNIKXrIN9aK0SlQF4D3Xhr/bRV797qWRJFcQr+mDkDg4Q
pY/udjlsWtdIRdB0tdE7G1AJ9j6JHYOdl5YazxqZqqqkZ/j8PpESM/P4JLXtXC+DlEpQd3xZEFHr
hPJUTmKqTsYM7wHRF8EbqBGl1+HBDO/hqL9S/pplnUJHwViO8SJtMQB3Tr8rG/gq5xgF+1mxkNCS
WN4bl8fHg5oGOJTLAomkaigYUpVxUs7Y44YMRxJacCGF1FwUpSE1TtzYsQJ2okCbOCPkAgsadK7F
j6+IPCcNBmdIDgeEcu3GViwNFBsTUhsUWV9lBa+a12U2uCm2LWB3JT/hVlHDRxA7Y+MGBMYQDjHV
xycRO5f0w+VHygKHlW7aCL69/rapTCuPgNwO7UtG4TStGnOpXvo2ZpUu3Zt/40WRihcDGsAHeon7
mVlk2/yQG9XiPfGTFTcigQ26lyTep5kHTmEa9b4PNEagToOp7fHlzCv3uL8xNUnaKf3sqIIb4EuM
C1aUYVsYSmGf0rBquUaGtwlCNLLOKL3vgzHWDknl4ALVGVW+DFA3P7s0GMsXHcSe1W8VDNHt3BRQ
GlEmkRGwl4CNV/DNNzXPDD515zhlcATtFyuqgQKX9ILaUi/uf/iVuiq6xrk5Bb+jiqIB0JuHtlA1
Qd2DLplcsF52kImyqKAi5gJVMmnSGGDZpMceVOcWSWGIjFzCzGTlr4gqkcIZ/5Okk2bf39lvVRZy
tfBccr+Z6xmNdBPHkDVq+VSC8c29KshLQSeUUw4kQp6axbyjvFscTMqyVPN6cz8IUyybMhVfms+h
lNAb7kRop/Jf8Crqg4Ba2nozB1gKdQuEpM0OGmiCbrB8IzaneJgMlbNZAlAhehkxHwyFiusnpvNB
4H7kkxjlsdPGqkiZnNGqBhD7bIZ8xoORrvR95nP/z5pa+MeL6AOX0yH+BiFum9QTdI5VJeuPOGWb
wm85FBtwOfBtWWUY8KFNP6BKQkGdVciTiQ9We4UWoYM3Q0ok6ZfeGHc1ChItG8/FahFN9ls2aEZE
Qp0CICqmF7X+2XjPArUsGcUoPh2tnobmxNjXMw8QVV/lRw/gGzEeFE25LQ9rWhNhJrRkSDW8sB/7
cPLpfvF1sUVUhFaVsoS1sPaTBoUiS2rOZdHDr+qxNUUBYp+8/HMXrVHTKDNyLtzbmscsbgyBWNOY
86jVMvRb16y4+QAUiDXxOOXV2hgcfLI19L9Wvx7wM5vbuHzatIO1nxfrIZMgB1fRr4tMYHmLFwFI
RXRoQHP49FEYnbD6x1n4ZMwP6SWA3ti0j4KlIpNkXmPdOIGrkFF1GupTo6Kk+VyL7VQoxSKovc6s
U7zvJ8VYqtFvBIMZna5bR/LWSD1h84+130oUHvVcgnzwB5LoMvdHkHyi7vRkVsV76ylq1l3eVvUk
XWwNLTtz3d3npwohRb8TOD4hp8K7klLPwemHOeEiH2+yOh/5vfPyPIuaLmLdwb5PWNZM9yNc42CN
Wy8FK7b7eC/jZczRgxx7W2nMTBADr8ByxR0LrwttPzncxJbguF4kfi9Pv9/RhkT6lVezibzb39pn
xOYWpvXjkjJUzu+/KV2ZHxXELcYeOOvod1KFRo7nLHJ5hlApIb4WahhXiS0Q3bDJ5PFe4Vo9dVdh
Vyc194mBEX8PRRKj/xQw0i/FVlMmiy9ZUuUlPLnu2bOylkDfnmbqfZ/EJW7uBhq+5650S5UO96f7
ZpEevabLQGeIYl0WQJ4wCB4V4d5pokEvscOCRMxZ1XzwGUsxlJ33uD9nxtVNNKAx+tMR0trzyIK2
WERGO5aKrwZyQv9xKXh0+KHW1VlyDNOGZUJ7BVfoupSXEwZo0JZUaemb09tPT4TLYpR2UCwlelan
c6gE/BKo4wGM3xHuPFjLZrlN8F0J33roMdCfe/JNP+SJoEWvpV0UxW3DlYihfwrFyyAx6Uu9xmu/
ujdAUbpJXahc5GoxWFZ/5h6NcIrW6bAbZvjHViAkaDnOWmUKbt3w4EWWcHlBS6TFo5rMemMG/l7G
l/MR/GmVofZ3JRhoWmr7h1L5NjSTMnRVadlbOPBbmB8XhBS84bOuiIbdzjOPru4Pa1JODriJQiDf
bI3nZOW31NIDFPRW0XJoWQ02b/sjmSZNyjdQVHVcuhbDN+WoKvthsoT2psfp7C0cGwZcuLVD3CIC
0/KS5MPg2Xr2Q93O3LCwSPWKfPUp4/pk4+t4lZVfCHW7fomt1uWtw68LcAD927EEot/+bCrBAM3o
58vCuYF5qh74SUGCpcU7mJHcyVXsr9WhCQDv60Kpd7p4QD/dgnczj5Yfl4J+Uc8otxHnkalC6JhU
ckpKXg2NiSP6zOLZWwP04zYzumatu89B+sVFpA2h3apn62BkHNCRl55XHH5JDlKd9rRN0a0jmteW
q26VpwYWGtDkJoGlhE1utKwmnLrbXvTB68/SozTwBt/3xZlrlqQ5ykcohFxcHx+fCWWi2Wyoy5aP
wxcRPCNdjLQtDPr0U0Uqx3ILh1WaG/62FjYhSvPEuK7aGptATTY6dcE/FLNMabWYaAdGk8wtdlG6
NmfDKtWWn3swCXbV/dYTzeZ0+fhysiyTXLQGAieuTLoaIqAePjMOVRIJrrEoZ4HWRbTzJ3sS0YhR
vyTR6m4C+x52JVGlSWNgUrKGGomHAHAr7rWqSjPt8EZShadWg7DQs/CQ2YhTUuNI7inWeeXkCryw
nAdT2co08gz7uw1TUj372QFB4I5eQ9pEKxkf6N2xElgnjovdkiKKCVxcSOvuoASNW0SGnMU2kkzz
hIncD8z8oDMX0hcQSQFWaL6pzy3Kzd3JYm5XipeEl74xjdnMFxhL+zl6iViT8wNj/CERYLdm9C60
obha2eSXVu8VkLrJNEufKAr2mPiCpz+Sx65ZMbJyalKwhIaBbv1Dr7oIbyGpLHozQKVlG3/Ls16f
VppFtZUaZo7RLTyn34wEknfwcW66zUzBHO9ygtVENzxxfgxubmMIGsvFGDN5AnJtMKjtLbJfOVgi
Q8wUrveZDjDMAqiRYsMlMcHToAKqmATLYE4esYi5hvTueeFtfQUBe+Z8gx/Di28kNKvoWLLibG0W
aLv845qT+0idFPAdIZxfl59iR3U+qS8xtn3qAe4DNZPa6BEnt/64YYW+zXK4fTInjvvRQSSV72Ab
pj7185uVNZ2uiKsbKMV1hkMhUx9v34pIWV5fZtyktoxYd5AVckqrq4cpFw/OZWePGdGIz1nmK3vL
/uFg+PmbXqxFwQ5TrOS8rJca6gZ/dN9c92wy3hcVAzKcA7DQ6nCpTRDi0BzzwxrIhNkVKw+YERNz
c+BZ7k4Glocsa+LVZdFgpfOtT2Ie47oD0/rIr/Y4FlaW/UwuyTIQIy9wBTXGsKa0M3i+TB17iQme
jlCtGNiIjce5AizJR7Ho2/Ajgy2waWsxpCLo7pIjnqJi72UyCsRpmWg9dVWWZXlF/wFd453jmIvB
QsY2dRYj9kK5A/ngvFGW5ftvuwyNkhQ/Jm4RMa/9do+urZxwocjC6a8BnQ//sHnkKaAhJpRAYj2t
bTJftHJp2VbU+E30il5eiIcuDGnQuNrxj2V4/OvNzQFwOo/mBPBzGbWl8X+ClyvPEuSwhKP+ENZE
s4zFb3k+Xkk0AhGLLXAkt0cvtOudpsPjEuaz/xKpN9UQdaK+SJFaYAVn4abpfqgwh2rqu/y2HNh1
2hGmp23nBpDjgWPXNqJd7U5PZWgnjeKrdsR0cy7ZbOHN3DBA6FJrGI7nlNjvUjkLx9aVyxVRWVq+
OAgcS30uV7DNXjow4JeT8PEwwhZ04UffeLXRKfIoqIqfJFfLKmh3ECUbmHbdS1QQdcnEbaJQGW9l
zTX0q1aQsOWroSp082OOwERXwVgIzAtOviLPxN7NcGCHPytd8GpentdU6WNRVe8H5OIvJQeyvuke
V8cZhSM+/GQ1xUhdlooJaD3M2gvMewgMwY2n3RaFtddbmvppAYrVOYWwppUqbrqt6phTj17id+52
zKp+ZPFucnx2O/D3O9khEhdNJvNdNcIVPSzGslvCAv+GBryFaqM6W9OHTUX9+v4doAsptacPG98j
1Q06Du5JBz8+Nz5IWn9hnEhrfUsyXsaijLo43ehzD+f1T14x4lO0LuLn0ZOB1XjMF5FWyeWeyy8g
g8x+vrAMPs+0WKUeGVw7Tf0kJkTJ7tiKmeUPrAjRZOrDGy08HEDls3DTDUlPbhEjvKJpE5wGilTW
SzoyqNScv94Wy+LuLf+qmYiAKnEIG+DQ4LAh8klaiux2+w3wRuRNCNERvPovOSgpbiHhZcOb3sb/
qlYKyebt31Tp67M4m+drcLpg3dztrj0UgLzk3uy4P+7FaABrFBQaMWUVQA09eAnNDFABWHd/mQMt
4rbP96jr/XLTd2c23Lm4LkO3r8WyDBvsTRuyohUEM++DkyIp9ds/Xfmene8WvojbGX45A33MLucB
L+wnTetmuE+JJnE/u3CdxBt2dAm40lUZs19lw+3ElCjJQGH9hNcj7a0SE31oYqw+1g8Hvr3gIG34
aUzCEQwVM/yJFFVWCqlmGezqUuD4Vbb0zbD3dH7zf5G7Lr6FJ+q1sDZrQKUhCCoRGMG1mc+Shfy4
14R6U+Zaf3+JMdjPh7UrzeaUopgEFUBFH7ozY07AQkFsDMTlpLQaweNhk0xQx9G1BDfzcPgiVUi1
A8LS+YEskSpiOEvW2ke6ghoHA74uiqR12mDiuJFuAECx7lgBUDYrgUufaU+RYnzG2+FLZTntEy4j
3w9/0L9UWovkjq0lOCzB/I1sero+ICl+Nx0VuPPHy/g5n5AFGUjfVEBi/prwW/vpqkC8+UetzeyB
OknlRSP6AVi1T4DWD1wLa7PUgZNCViDpQDWA736LFkhTfI5siSIAjFHNmrq4NT1KP8JKKPYOmciV
SThPS34Q4bKmIRUuGyS6+MuZ6ekOzAHj3LEwNWGyliOCT3UsfKD1/qG/Zom0rY6p6Ea60XLNDXy8
HuBlIlFBHl2Bzsb2csTo6v5+RpviEAabSqWkkHI4+2e8k5z9YJ6Ni7s0PfjWuARZNsu67w+gZ7lb
ujsKpSothAa72n1zt1nVSyvid0Lp55zeVyuBLurPpexUgPv9eS0Vv6FM55zo3VX15j/XQdKv4Hbt
XQLbpS1PRCCookeB/8QB3doU8r3sngNweDjbR80da27TW6QowHT8KisUkd9LGOWpb+WNcJr3Oj/l
jYoJEU5Nv10PMJPNJB2Yb0Zulm1qUA4qNpiNEXvWvlCMI/VN9wJzPs2LV5KuNpclvDc0mKeIQ/PH
rFMnOigqE0lGv7vfyugNygOCPmrAc0UhXaP8IrtFoT3P9zwROypR6atZe2sPk8ms5h2JRmKvYf8b
PLbqOHrjjRwJYTgGkmkCntLzlYqbDhwadUa71rBg1KDE359XQeFyw+Hc+sWP2vFxXG8CzEwSDDt9
6QWHRdMkOv6yxTAMRNXu0QB3kPk6i3CA+hdyGrl6UvWGZIlmiFcRCoQEmPb7nV7+RopBpp7RiIaB
5qXt+iJPprbzh7hI/B+mi8dsb63JGrCW0NuP4y38+P9k1+IDX+lhPaOMRvdgiPKtOORhKZ6SVQqc
tG5G4642j1D0jAGuxT1J9QoXk4prUmkOYVVZusepDXijyOP6mH8nXy8wF7JKGuk4+pCaji+jWshc
vT6fmJ+K7PTtMN3U+aKBM1S08Js/7+mA2wciYDZhHFHnECNq9fzZhYwA16A5FaempxxKpaPVYdqT
5na0rEIW0mSyUcoqzXb40wQVCOok77foXgxMczmHNjfAZBl7X/oMgZdtZGjEm3H58sDjAW0mTFXG
+E/wI0iVE+Z9xW12V2tR2XHNt0j/wne7MWGIWURMawfP645XDCFsQ2pC82qJhEAckz5l84zAqwzj
tvQ3eVR2E2r63IvwCs0XQ8aBrjDeEVTxZcNrtnFo9U8eGJIFG8TDh+C96K+Mt+hYsnTjoM41Ueoo
J1Oa9OYuGM83JkHRtTN5QVqbkMi8VJ9GWsoQ3e6+m9ur3C8gMrjjpJPDY8gzbZrAeZ+OowpdJjEJ
v8AO8rwDsF0TKwyWpeb4Nu4JGu4XurgM8fP9FwVF7xg7dgDolYy0817SjJzHAxH5ZB6cTbkDMX3a
QxtjXeBkgo+MG5R5fG8blWp2fznUuVWJ/MJY5VSHJi1213932I4HYFucPfkah2WgSPCSudHWlWJj
w2kDG3YVyX+PYp20S7ES/LPNIeznQtqw6Tibaka2AbyOVO5Wj8fikhdEtC7fbfSB2XFSoPqlgkTP
k5ZxVIQTgvSfgWo0/96ggKnSEmU1XHcK0PhW2pmTvZyqKL47K7eVgmGZBb+eRi+GljAsquh7ieQq
cAsTdyCgNYK7GVi58BU2GgOHdHZACAt50rDVusVVYK7w9KHGd/QdQoA/qTnrdsKcbdGDgXcpFHy+
v0lazGXJDX0ENPIIr7eb1vjbr86tR8lO2neQJV+5ZzHcQ5IT8qo2v1ifExlLc3wNYqlmlfqp1eqj
NK7KNHaYvxjDPrWW/sg/W2jc+TYhBuUJls+4LDH/gkZAOuO7gw67wpR0aWa9QxIaXa4eZ7xhjx0P
sAEPPd6A2AGAdSqAm6bF1Otkofxo01EvvT0dTx7EjIBQeuRsCLwK+g42yQnBLi45pwbUfO5bcIth
BGiOws/Q/0YqY9RuCOPkgafkyPULsPCCzVhI0pIHSrERo8JhOdhPK5bJnc5LIAy5RohtZdxpCDpG
b/ibzWWzezm3Myc+YS7JEpxK1m4rECUsaujZeDlwFg5XWLx7Fq5YaoMsgC7tLJEbhNvZXa3kZ6is
nZ2Q+sWu17hjFaAHRsReTOijdvcfGtSAUICBl2hLNib5y1V/q7URmfSC1FJWVdaRRAE9PEsL+6TZ
v6XSY2RJfMm98SmbHCsw4YhBbctB6zntQ1ITJXboGGouXZmLGK2UgsPzEBa4K1VCeBJzdAyoICPZ
8CwJ6cDgTDk89uWfli3aYPZJ+8qZTXT+yYTSwZqyxFFAe22l94aEkciq3077SRPbYitRUgHZWK0p
qQd+CNVjCQXD0L6MyJN8Qd+dBTvXIJFEox2KqzgDjhtNjaq0TLKPXjZVHdiqgGqiZcOKxPAkijnq
jITbRPWqMJGLXrWqti+wpORLvcUIDaAOaSmReTws/Xt4gGoqr3qFn5h1+mj++w/H0DZOikrEBd2v
oOU6E67Yw895hISd/TsZiqcybvbBcU6NoG14iMZaoX7B1bbTjiymoG3osYbM3whA086DeIcPQKI6
d9GCDalW0RZmePsujHD6pVF7Kt7cnLkGNhkIh4aWvvrVjR3K4st5ZhKvlusx0LowxNSeo0uanAbw
O0wObZLuHfou2zHXNewhuMsa7oixkDb5isYGXpLZxIQZVVHXzuzDbxZkqFyitF6JFfYH3hHZ6seg
r8Knep6MtBniiAc0Q2ISfbe0JGPkSOcUyMAh4oXOt6jDZLK7RiaPcTDbxZ7rgVa7fkYSIAYV5D6x
BlRKbwpH6iZjoxHm1USScb9kVUl3fj9GRF7abas1GhJzwxl2moU7qmIfCgPOOkFpJkgMXc3qlVZT
w05rvEI9dgYngyv6JOFVIpvFVjafrekuVHRMv+zQVkJwAiHcX7uhiMHg4MbywoKJvvZdDSfoxXWp
+eRGWIsMcsBdtBZRaoRhJ2zY8doTy2//7ws4kOpHc9io5lAM/Iregk8wQldELgfnKJWdIYut2TDM
rVkT0PncQm99Jj5mD1VHKDN8tHZzDqVXu94csGmUi4sbuM8jIVoz38zDHrzdrK2D/9R9Ji6ssNFQ
nxvXPmcmIhjo4d2u4wfxDBkcXxmKKqAkk2cshuxD227S29bENIiA96GRMsXtVXOTDD9Fgkzm/unA
/E8NHJIcPQSb/dqYogwCu2D9HO8w2fXT7ppj/qZXYknZX+yZr05lRLaJLmcbsusbQFq6ol/lqosz
4geJOrAMhXjUIWlNLzMR4CzHLx8TmTDRw6V51sl5MN1Q6aXjqnnVkJC1jzRKKmJGyAwBaiw2PFCg
isABzdAutNr9eWBzZ1KRub0YjCGjWqpiZzfuJdxx64wQCD+EVSpeSkhvccp4tCfjZYc77TrxZVQS
ro1XpeN27YzksXhWOrc3o5+IW5Jn7A2Ed+SMcTLC+JB3LzojiyJCpSWse+keZJpgKGLDo/X9eDA0
G0kuTa4FV7qjiG5UCSvjzTvqDxFxIVUIJez9lcszy+4aXCHFk26ZMo6Azm5/LQiY8EEdngM8iCyK
MXpF6a27/Aiu6o25XffhuN9Fu7ToZq6r2Ggz5ttyoIRJ14DB3yjSFyjMld1wIFu1uQpNrdrZi2Qu
/gsi3mgQqFjvQ4VON+N0b/gSqeCj0jTrxUSk6PWFxRur6sKTgUOmUCYIxQ39PBEPWu/+D90dNDRC
lHNaZHySsAi6vDj8atuhSnABgm5PSYvs8ojL9W6v/sh4QH0cj6H6aLtTA31dlLEBbj+LtSwYsivd
VeLEhQNYRn7MiqzoHnZsuVvhgiuf9i+v8xRFvT3xn9K5kNKqxh2+AZ7AROdAaQ5GNTEv/YoVERKQ
jSR3slxa7g6KyqcrfIDBCOf0RMyFdhBubHJRQ/6ulMPWCKOxKDL27qZHEzn7vSKHbZgCAtm723vi
fNV3iAYc3h+I6LiRnMiahWMA0S3fgOFoOC83zlJ+X3gaUeHLufg4rNEFoZMlUDGWHJM7JoLreNRg
f0UjB43jyspii/IisuXRwdIDR6C5bDK3bvKSgOBKmWBDm+7WZztcc+s3YT1B2c5C5/d8RlWA+jcc
g6TF8rkoYce/e4s3EBTC2SccDwxb+u8ZpwzlCyW3OWC4gAl8MnV2KcAcGWlMiGoFjFqi4bAAB+0O
a36Apst1rAjHqO1tmC3tz7Da8rKQbH1ecJkae5FPla+iR79YR5jp/aR89r7L6VwpUov+twXsAKEr
MKxGmQl8awlK0vV5h9SO9jReZrFB6dFiDKNHiW0sdkckcCC/JH6SY8rgqRHfUzYgpGmIQ5pzMckv
CMeAbR/hcW7PxxMIUQ/Hu/Na1uVs8Z4ScLDHSrsAZWyaV+yQjXxjec4U+SMjgw3VbUBxxnCma89s
PX3t3jsIXsNlNd6lvPwIsv+e+XXnhS7t2xsGjQe7m2IJ/uyJZgmbiF+raiGsyUgRB/6a5c6sV1+A
dP3hxPGM8UuvMTNL/Mn05RreYmOfOhmkBJLgv/Fy4SgC9lWfc7+D1vdDpeh7t9B2O41Zae6QmmfL
sw2W/TrJob8KNgfgFqaYYtf/n9RU3mgO1rmNs9G0qw6HRXtA9nSjRgTPbVLX6o0ulyR+j9FZCN+D
R3wA9f3++anLSHTs0LF7uHS07KMk6iHXVJx0+lppBozgCffhUOnDbgSi/CRLxG8e5wqh0UjED3zW
w0WTKm9PChinZnWHAIaH25PNTejRxw4fLkvj1ffpt1Qvk5ZOFnb+zbZSETXPZIqUsMhBVGuwOriY
5rCNdrWUkW+WAp2/dwnCs2p31l9g6KTrAWTwtFxnQ43TgsnJY4OBZn7dijavXo6ASEJIViCzEBWf
X3ZOFGZjyoC1Fn1Vq1EB/VgqgFmha9EwdXvcBUPEx/eWkfb07jzLuU1PB3NbRuOTLjJDfaD5JP1W
eUsv+CIyZ2of0Y77u3b3YL8ZlGzIXjvR0OHkWEQzoyQrB90d9DsRcMPOmS/h/OTFzLjPE1BMTg/3
vPrYtQmcnrtpGrEgXhsHqx5BWDRvgQLBzUzxUd3pk3hdlYFPjWM4t3O1LLHrNn/8SLWAX0LC8N4G
HM80cEKFFl8udj8TOaSTtaENZso9eKn+0WJcpPwHflNAYLPQIQr5Tkx3e3Wt/y5KmVnsEAfbskIo
1HOiOWswdMVFdkepry0bHSpcKYIoqhO0ocbxWejUuZ+3hax9eH8gRwsL+p5lBjtFhdJos/I5663L
8dShlC6Tx4SlrBymDepCGRsJCFAU+UAE7Ap59w724EdkRLqLjYIH4GAYmEZisdQ7Vdeaw+EKHiMM
s5XWb6+PbLZw1MZz7/hSv2Zt79UikyIVc+Y0gmKglVNHhGTq1rjAE/T/SfTuukgvLnTbd4uGECT/
G+bI08dHIXMD0EOYWPyZzmlKZeabmQAKZcrsUF2ECa7mpFV/LQ3RtBXQrO8p0aKS6+PNsXjwEtiJ
xZ6baTZQwC1Fvbr+mRTj5ewWeeI2mk50tZKf2110soS3iDJzZLL9UflJbp950RTYqcwPrPhs6gsB
btpM+EluEUUh5NFCoB7YP8zjGw1t0IE6MhbzjXYrwE2adC/1LGjHHxJVxqb9KK0szx1E45fYGcGY
TfrZr5RjMqrouKrZAzmXtUGtUJgASSJ+NTqua7Lji6UwY3bi1p6rsUwzU+JzIJ0xXJiiLMsS86P+
FSzt1jrie3TZzsf/klbfU2pHFBTjJfdZrNZRUeyMWtcjwCXvaTX+KTD+hhqa5E8bB6lu2Zwm+1Kb
OuA/mZ3vUiNZ2z3ypTb7ia7iY1h28e2LPt/1eUQExsYfoCJRtfNUFtbpZbmh3mhfQjawfZC1t+ll
oebQMqUWm7W8aurpczvi543uK2Eysp9q7CIxKyYwbq72sSNwCmxvMJjFP6rSQdSVSqwEWxbof6qf
ckmCP1SDK3StVSWqsE+LnkpL3IC20Vuhe+u/NdjVu0Z/rH6CZ2TSc61OGqmhYoVko7g5gySDWflB
L7ESFfKXab2NnbUjq4fmnvpqTEFW4pMGOjpaBPdnZ6f/I0LOFlQLupvnj5MCWitOKZss8yE/lnu/
dt5Q0hVj6jLYK1co9mAkOxHjYkgNhvzCNJKTm3rmGlRHlK8+GcKNdwaSzmPKpIzxg5MaMF888MMS
6uyl1E3TH+nJXyu+HztyiAWGamvoyQwdAkAtAt5Qnank/bJ0olHAsEW4bupmTy/lvWmHg3eLzWNS
n06kuZuDOU+Od4Cm1WW4/EAlp4hqs8fsJpbxHwzbVCW3arzImS2e0eq0wkzUFXu32WfWQe9N74Rq
rSU/eSM8BbKSXbfbxAl2c6yNo9EeCvZgebCbWQXFPfg9/CgFmBpwK/mQ/46CfYRIzA2hooJUnoZf
xozFrIM8wSPuo4/9+FykMiR73y3YQJ27Ye/lI87RMZdsZguDYDWaooaOQFffvCJXEgLgwoeAeqJb
xlPV8+l3jUX+uPnOETFP1Y89X1akDcqLjZh3mNdraKIXEsJ9vgsBkU7we5clFuAZgoq6ruUqCXPS
VQKKrcij0FD8hN+Gcv3gPnv3Td2gifTnUl589X83IAFZvo43xNcG5mMcsaHH/jV1g4nZTMgYwdmE
gSkGKDLctqCz38JE6Ckk4yvhXXXGf+6t0evmFMp1n/2MJkHnYYu8T7mYQh4kfkajVNshppeN5UHn
XmaB62CGq77bL7obOXY2EyPsJSJ3M7CRj95eZ5Syb9UgTeSwPxUTiOdnA4VbeHND7UXs4OIrSWzT
g0/vSBFLEqL8TXQ5LZG2Y5l9H2oxkz0WgHU/kf7QxlZgUtM+bSNhJfTdgxxnO6xQMvNtk/jFJZBw
ihEYMTI9Q+mZvC1zvhKkzBjHh+HxNdNfL5RXb54sOBZB0gvELLx0VnuCZawUCAwFa7eA1SLZ5CJt
Lop9hwVkF+3U5S3+q0kvmPEUpWDzpvuQfQ+CUuuPu/XU5AEDPu2AUpwOHxfpXsa1qWHLGU67J6NW
/9TARA9sC/WUJR1wAOeTpHJ9qZ7jbx68wNVzDER/ZFg88sgzfvjLQiPosKi5duoK3A+srzTZtT7y
5/rSDd35Jlsd390/WfjpLXo7bgaGY/UsMjJEvW+gmylI+xZ61cv0pf9NjZM0QCVeDorbSSNOuABu
/4uM49fvhQX6GDfwkBehjS+16PY9cmSU+Ap3hoCFrvZFx3NDq7+PsaOAM5nQ/Yyj7sb01KSKRuR4
1q8LS9C0jFJmA3PL88PIOxNaHdu3YFhVoM50B8BfTNiRqWbwngGThHFwnr6jh2CJnr7A1HjqZApj
lRXXc1RoqQn1sPKkyM/7QnAFvjjqTY9prbyqVwZeqLqZoz4efQmiAWifwxNfz+SXcUwKVB6n+yho
o8ouB2uy4FdpdpiIEHwA4+d4aOO/yOTdONEstX0bvKuFf4zLEmVBDr/eYCaGTQPBVyg7qxZhYdd2
m9SbAFKSb/J7wwrNedaJTcStosDhrBQ5MRpkdayypJR2atGPbIStz9TtOy8PnLQxFwaNJvjf+Ibb
ZzNxbaegLqdTE+85kQ9vZZ79z2JQJptEupiUe2vYEdjhkN9+M4qVv829HDk/+tGrYqSt1588csTx
+BMwGYh7sHov3bNFChEJfJAvWWX7JvCeaCMZIRBX/D6gWMD9l5DT/kKg6h2ZeVextGWUNIg5tiCG
1nkF3QKXJDHitOwzW3bER3KLiJPKqzS/qBX7MxwQ+p0snTycr66vBTF3XwShq/nRy4mR6vEm2LOr
j6AU2S1YDIy5aCgQLdyuT1mqEQkYjdsCHOe9CCl+BYob+fY7yd6pqluAauyYbzahVpShVdMXTwgS
ebQE8maVReyBvGSTvrsHgS+u60Rm7kR4xltOk5n7eW2ELenEWx9KiDm2VOCAHGDpIPZl+kRnPA+c
ZG/WhdqWKnrTdHEQ4A4wKAvuS+bew27/uhH9OumM9x1xwwBdqv/EkP07P4UJZZBy4ZERcGkWAalt
l/K6WHhhDkiaoK8neQDzMGfiL1vAsg51DiuL4vRFrDXGZnpPAKp4bVjkwjIn7XRQ2Za7dttp8BV1
+QvlZcJf61GGrrZCNKpMSP/0IbfSVQUfcwVN2gUQakgiBOwHV1O+fUp1FnYWovojEwz6Z00rItDx
fPC3yVSvp2WWt9v77DDoN33B8I4K3Ks3iMh8Btb/xRdHb7EmV94rzNXqxokPUMF2mV4ZIPP+IWLx
aFHTgFRd7Vooo1VXapVWAyhJvjZoWUnVUposXUEhGfJlBK9a1615rAmLaiuGUBWPbEEfNxLt2YBP
FZr8GbN5HV8UBXjfVk0cnrQ7t2yW1/ohpiKm9wKNwG9KfuKMoFCzvQn9PlAtdebSiMmQBHPQvCCq
fwblWa3J2D7ImyemqRQDX1eD8tOr7WJ0lf4Lbmp21vA9umUWOvmSS51RwDrD8zHelYcab4Hdw/Rt
GvOMkBcnTupJLtdYx6MPZ/H1KT8menSC9qYTFnv/h+y+357NCirdLx/pntZ4HYYMNTou8Pd46yN+
6bg9UZie3ngzf5rFRnzELiF7EEnC2nsIWQYxJkynOoHCOSNdovaLcHhc+vf5fbxTliao5P4MkHqI
DLQT86VyHce/Y9pGcaj9L+0hg6KOektSaYD76hBGPHXYL+dETK8zyjixnjjpbtnqIJS+kF/Y/wKb
UxXW1kl3f1n7w/2ZVsDdr23l6xK1fIKugr0WS6k+aP652Uepz2z15SspcN4Zz5eQd7vv5BzKO3eq
fJ7B0EPB8LnSJijJyt3UTRlX9YVUQ45aaMjr6VVAwGwVFAwSRfUFF0IRIaRLQvPfDjz6bNXg0hDY
3iyPBRzhS79X3JKVcIbwrn+QSezs8HUmYUxIjNsd91RqDPMqh88v5oJYuwO5IrG8l+i+ZZYyaqHz
+BI7Wov3PToJIKOovmphe+ULJloNAhzzSB5uwKFF4dvKGg+YaULNDEFnD/N6tMPLluhO2Nn5Jbd2
lmu1kZspAJ1csTAxloGXLRWXHwIV45evn6AIwW6Q7XYoDx/l69jvgr3vZha2zx83cMsaOU1ZripR
FGjOsvthQc3axKOxhoLDoubltwSb5gfmKQnUq6CtsTmsl3WkTUMmYAi/b7UEaTvuOzxlVMBIEYlA
Iw12HDo7xJ6HAJ5aYnCUn7Hjks49sNA/tYm+KWijdVIctxvU1PjfTvl+628oKXGuUk6lOi/gfpEA
LRxcPx5jcd/6sGUvOT4k/gqxqbRhlnE6HtS+oKJ/wuB/RY4M+cd3R1lk2SPIMRsyXKW24Q/3Do1r
dUPhB+QIM631wp+zfLVxcvYJWNYma3szA0HbayS7E3IeALu5H421INiX1fGPUe3ES1MloUjg4Ay8
LdosDTWQq0UOmULJ8ezmI57HY5nnSgBOgd0qGjdG4Bu/QZ558B0jS1L0QlIh1vE9ZCOqDTHt11B9
rX0+X7ROjw2PBZNgOdvQgMmnonKphnpweJKRORLLEe7JIqQI6tVVsGi/2u1Trs23GDQCVMiYNOSW
KWwStKL1IOvJtzf7/0h9KVt7L2Vv3GdKHk+tb8P8Glbqoipwl2K1C10DtcdNqqSV/G4LX4h5KSIt
drXzzzA9+5Nis5wLRjWFUGoCSmZMTKQE9cZNkEWMEjOKiNkslNYFDLm+d1u34xACWcsOSM88dKsn
ogAn8JvJKP3IyU/35qtv1I3foUciy3QfHv1dmOd4bWtNm5cna+QIv625xP441ZnwHwf2mueaa6Qi
IkDwnk4Qe0Rr2akqpGGTuRXyiD4K8bGb3xaZcmsKdoWPSCQ7IF9mrnmu0SrOdnZOCObe+vZUpruN
xx07JJ1HjsP5EKD40GArxIhCccKLfon2CnjmU6A9U7NmJrHKa7DmTSsVIKn2BFE8U/BhXXMcYlV6
lMNogUKQqvkWIwF/hkAAZIwJ4ksET9lw6pGdTRF7M1rUZ5OBSQSBRp6CdagMJzyPsWTEd04IMcqa
xXNRv600h9kcPHHj+RX2X5L/hCECXsHPBOwLAyOaqdjXn7fHEHTNwhWDfZgz/TyZFKcY4EtmeUVt
fr9V3JPW0+tEjumD7D1lLuYTlATCPHvwy06Rt8BHmi9nLE4sB21EjEJPBU3XRu570SA3sZr166A/
UGr5bobAFiAYSg1y61KsnmBBLsxa/PbQXq9cGaxkrMewInPdpzdv0WAjZviail+I4CMKYcy1lOno
9rdbHWxJJuqkpcxjhQkhOBCRNMdbJtVWx3bQs3Fct9ol5Yx54gfMASD2jr99o8PntkWD2k78CkCs
FhIBMhG85PL10qZl/ClCBgcK9JsZCrtmIAQTjripVSoka2+4rdIx8H9TAZov3CM1yzm4sg97/FUu
JY+FEIEfnSVrdOPa+UNGk/dxHDUfyquwoHdhcqgBr+ehNONhB3CpfbBy/9ett2nRM1J5YKoWNNQH
tQr4CbJHO72EZOJVFok3RjlrAXiQi3Xezj/buWgTBmMH4ZsGvIGqLQmS9WKwnE4n/MN6+Ootm6MB
Q8dRe0soxNWfy0p3pBzprWG+IyDMhmgm2omzoArv0wx22hKv1GvqHTZ4+Vo7jvl5kgvHzoQpN7rG
hGdIWLRczjDk+ncsYT6DIaHm9ms8cXf8VdWNTLB4g1oKEVwMB6dOIrQag5KWS1k5JOsu/6woDeCV
LCk9zn0KP6/Y8eb68D+2xRl+acOyr9CoWFYv7mcJKRT5mxx52/Lm/RgA9f6l/xn+G27ix2YlYFn+
Lg1a4ewDnns0uJltrrv/b7RISY2vg56w9G/16YEt1kc2hUiPfs5NiUU7Ui+QjM8ElLGjJBkWdPW5
qQULB2cHcewXyLNelzjgmGr1ZdSOCZaAHLJKnlTyAq+ndr1i6t9zjMHTkjrVA/o4pcPQc47/hPAX
KDohJVDMpOFww2EZQFobd8A5nwG/ERnGsqp1nJFF52ogajNjUAOEMXmXJHKBpoEdReIy5ccPI1CS
4KuFOT+30YRJ3qfjeJjmYXP7I+zr4S9SH0CpOgyw/l/m2F2MpF4bFAwqH7Svw4bdaEc/gBAJ8zmZ
ILoJYE7ui6qG2zp8Ruzs/5zDMye+EkClITV8h7mLqts/xCpYNWOdUAvU9Y1ALUkLzQpCCh7YZhGS
GeE56acsJuZUmgfTnXxf4vjLCAoVksabgUtShLwJviWpDxGzp+ftmvz3nxwOpMM87FOaraU9N/o6
6960f44Dv1uooXZvoam7hnL7PS0LPIWi7zsm//MpLJF8UoL+ivOVJ3kWux8N3QtWPshSxTE83G/E
UG6MnZLsTQHSzj+Lgwvm1/pePwFnpFyB/JZ2Ey7l6trEU3iBf/aETlRnVayI0FW6UnIb6EgVyX2V
DMj0Ibm4aPy5lyqfHwwu5uPoQ7RV0aSR1oepcA2Xc3RPEGl30S/mRio0LTHEl8SJ8t2E0fYbNUFe
HqpiBEl8LZbFFUZ3Bs/Zsv2WpyXA6JVAnlHJd49SotQTtJzu/tkOw+Jvj1FLUCoE94H7+I5Oyest
i0FATCKhwlIefAsovwhkSBVF4tadGzP61zyQGm4muUH4iZswl9urWMHh3/ubCOFRxWKjtbiiames
Ji+nAGuHFPi1MVYaYx1yfGTcMFpzDx0MN3IZcmnkiWsTP6ORlb743eatJFce1qaqXrGiNYiUBml5
KWyzgwlHIrmRpCOCxPDmPDFcrE0AR1D18Ri02g7MDB835D2w+C1KEsEjF7kcczNzXWy/RSn0dRcZ
6ZSnlr/oJRUSbbErVY65g7x9xyvnxiYP/59DiSRnPkkDqHYr6CYzakwUnVZCiZPj4k8RiZnYZE/B
iOUN75ug48WneJutF017wI5d5olo/4Xz//UHyie5A+fRYsPCePannkJKPz/u8CMQxF23USs64NcX
MFIE7xjNaYwiFfoQ52aqMsGYJgT2MZP3oTJXd+jZ1GYDRPUJysr8wIJnBAUpq+1Fsx7ors+PwAqf
/KBCNeNYKgROmSH16vwBY+NbB25ZBfsEBihcf7LMFTsA4pNBgPLU596gRSpSyvs2LWaCi8oCQleZ
Ns1ZsRpw2KpXU5BeLJAVGO+l1PgVZdUi/4+XjgR8v6psWgtcI/UCloyzpiMWXTRqNtKcC7gXiprF
4ZQLQvaSWPBVMi6/M17K5PYBqug9Rgz71YxVzrC74evrsHcM9FyZ8HFdrFIchB7tg/ZW1WAPDC6e
6v3xbTgYrti4Oo8LBJg4gRI5ggFpIOSyOY2J2lYbQ/hctFvxW0rOqW8vpI5dhc3YJCdEw30vTwD0
8hkaGl8+24w2QBwYMLCrcmakOQyW6YJV6+KWn0zMaV7tMdliVP4x3YN/Hxw/zopFrwXqBC1uEaeJ
Pm2zhmtg9pYrjPkEkUviQG+c86jcHysH350hhfj6jD7sBDe/aNN7CXLcxc8u9cn6AnTuH6lTsABo
WLPtjv34jsGt9ybsxQpPaADEcXa04tH0Tv5S9ZnbHJ3lL2OkSNgDBaBCgFFk5isItWnj/bnMbBbg
eX2e4XxJHYJjJiOqhrl6UkXs080IAeX4mHFfiJLTYlnzevsZMjV2sLiTNgXj6mmue975RCZV/Tdm
Uhy77V4cnQ3HH1WC6dPtjP8rrvNQzI3VViisnvXCR45ZVYgmWpIeh38fBq5BdNsHU6WfU21uS6cH
z40X6w/DZqDiBYWwZnG6Kb3cr551qgTja0KvDwjciVLvyh5L0d/y8TO071X0Y0+nX/XW+TlPXH5H
5I5Y+04irLr2g+E5rjrzOGfAJcOTwOVwzU2JUR83LulUXShHSLvmfpzBWwdsloSN+/mcV6Smgulk
qIfZYVIJc7gZKOv1GdV3etaIjF1UvpC2f9qDjKnXgTaEwesadezeBil0wTuvBHQSSb21lRAPOyuT
oHTapxBa8y+O3L+1KR1rsz+QJmbWPpfNH4IwDUrL67sSDDPo5YrNDRz6DC/LTo2ZDBifDQqmLENa
LCPVEhd1CorrWaX6tPn684xOlf3KBdwZHdvW9U77TPuWW4JlkUVpCSV4cb0Y7V7/OMTe90rFwNDN
s+4b+vNZRvS29PgVMo6KvzO+LwY+e/cTEiug5rNqISFgNWc92Ow62mB/rsBv6MgVS6ViJfhfxyZD
2Yv961GxZhB4lYCAVzqnWSVfRiMc2VJaiIPKuZT0ys0c2UXU7Sk55H9p2DcXVPzY0qhwC9aPIBO3
GwS4+iOQIk6mXkbX6E4NSLaTKu2hqc9y8QhhnMyioIMQyxbnTpzUegX6HYVyJ/vV97XsFyXsn3Mx
87AnyIhMcCknSbLHnpO4H4f+2JXt+lmm0JU4kI4hTAlnAxyNzFgmMgFPCFWwMZFZkXAW6pTJX1Zw
vIFymqAVrRSz5Ji0ysfhAj60H9giLPiBOU62bxly/iU8kjm33gemCOJpZd2vGIL9xoo2oQFVincr
U7244JTIv3Egf5ncf0ooRDzUwsRGZIM+0H1+EaL8y6lxbkOrEKgyiblnora420ySOlsvLaQKTWqG
I6jiCpOpKO36f3oEyzXxyNK0VejDixGrV/t7fuidYcNEO2RH3bL7LsPz396fDVWCaVrw7gRoWzyr
RWjaYHYxFYJuZfn9mI93MlzFtAWlcwi7HquI0DDWbiPOkhjeh/pHEmd5w7197iNkSZwzloxVZnrp
rvXsv1iegThdYOI/EEExmlmYb99hEW2gRZrmaQZVTDZ1/G6KPF7AhBH0NwauKLH47gRb/nXQhn/M
AqAtUYdsVCQ+NiTmcJgxzYpd3Pj2bAoEQraNgro1HGcD/tvtSFMjzXdr2aL2Bg58W8FHGR1Rxt6T
zoidudq54amgTBqEb8o39Ys821cVhLYQ+dnw/qKOl9uSVzgsIc7XLBfiqubn5KTyI+xmLw68dXRN
VSE3xMDmbvbNLcN9qxh984eXyohxpFKRoBD2rjSQJsshdy0SN+9a7fMgt3dRc2vOXzwnxjTiv4uw
+htw5ewrCxFmOzDl1chv0iLaAdgFRXJrDsakY/GYfPTqUd8LHVQ0W1vR63V87nLeLXgMZ2glaXmx
8PfmMPx5IgS0vfPlse9Vp/W+JTPzrGLW/ByiiunpNzwFc6ouCrOX51KhmQ2l0fT15hj4/GYf0N/R
NXGybwCpEMTIlFlVsu9pHtNalJIcYbuyJacGQdOQeYk1i0nR1cSSwcP+DpPFMfS7FuM6Pjq2X3Pa
nDdfsSG+RLUi8O7KqD/671gBIKeISKN0UZIA4KA4J9wUGS0uKmnfovNuQfHrfk+dCd5XVlbLaywi
Dz2d9aAwUraIATdM/yb58Mx4lKCWhSmTlgZLr+hbrmETmruU+vxvb1VGsv4EZt8rCJDzN1ukDMjG
WXQGTtySBxfdre682yHKrMxy2LQJJggQVfCrghw2IeAZmV/EsomtObfWDarEPDiQMv0IbXVIc1cU
gXkAopr0wZ5s0d+VZFZsKevbHpadkcm1sMHeOQqwjJZCQRYD20d8Yepctn93gXw6Wc0liS/8yN3N
A8lPu7a0QfRK6+3iyK0k0ZrnuzhuwKHjC1jvHeEyNpdjFQ0AVYNkj0kY+fh1dPvj/DEREezbsTNU
IGiNql62iuPTuRbRe1tJxAXREBO557VYzaYJI1RyJJjPwk+sgyBGvFc/mXx1Eqk6mxB4Rrpcd50+
uwBsplaa+mvwxakJeJ6EpSg7qGRwpyuuVDABVkBsjVRaOu1Wl/Ttmqp+z6aNTwZBvfQOJ3vNkCFi
zQelJYn/8/WBRcPpP4oeCt7TTD+H+90cyPvj8tZawO2KONpnRcLWyw+g4BK3Spv6ABO7cEBI0ymU
ywoaLLNNIKPTedQ77L4Z/rLalzUvQIkYx7W1GfiW0ymaQAvzCKxSfvMua48pJrxqLzR8zSQYmm5F
3+uRNcSkedLg9r0+wO5LvEjqYbmOVeEnQdgALrqxCBcFuAQD28+NiymUhr6GIZI0OkwDgYoXKa6f
Xyww+e4zEJBZVYoIOlNu8Xpgc0gSwghMmpAdDPzbDaFFum3OEaAkgrUhsNA4+dK6AkHoxEPxajnh
wXrcCHmh4u+haGtjVyjOUNn9PQYoxfqsvjNwyCOz5khVB35b2+16CDLDd5sVFmOFiVOrY6ttHl6/
SwhINDKn+LFICzDCCBv2k0YOFu46buN42fvAfzuWiKGMPDO8/3/JTSph/z28an7scSRNSHSVTGem
JnAAR6qC/2TwO4EJ6oKGGFGa3NEPryBeIU8OATuX/hjrdly6soIYHqfsjsKiieNOvhYiI2vYzSvw
xqyk/bHTsne2fnzx7aXxyXtADXML7r1t7A4E/eZSdBHFNEAJ0GrKFnr/90RyG5HyCWZS8POFWe7k
uZuy47r2/RC9jtCJRKuX6z4a1A9oq38H5K7xQHhcvFuO7FSStyWWyXGAxBxfCxqDZI8T3YOp6kGk
cbxTZ4Nwf60HElUIOSeZVvVYB6oFgDkCgXjvHvMzV9VE5XccOx2d0pIpm9cvy3R2/9Ik5SDNlbNN
iLVMA3/mizwtGNZGK0w3sGf4xt/R/eOZgimkCCSbXMk9uGOayAnGAeHig8oc9lFr50fLNPvKWAC4
zzfmLsYlPZvfYsanHFyeNuYkNxtBqWTN+YBprwFTMANsz1jxiWWfvnRL4RHa6vBuonljD1IR0NAX
Vm8bVEDI7Sm2sxtk0An/khepnCNQuQqWU+aPbVgFtQgErZxVFSCUPG3FCTZQJegppezuyqz9trMD
L1xiuojM1KRMLD07RlFrLxbnCHB7t/OXt3vmU2vX45ys6tMYSch9h0A7XkrVgl2WnygOy/K1Xv1q
u5EQO++zOtZIjyKUbnXxkthI9RQu5cRs0N2JT2js+OVe1YzTW1JU42pY+pdKz6ZxJ94zo62JJwiE
r6GJPdL5DjOk1q7AonHA2Hg6Ky0xvEb0fSuavqYTX6ZJLdWq1/qDomNW+d8yKg0YdRgc8X7pSGZn
etoohNzz7EJF67yFRo/6Sc4eCXlNytRswaS/EIToGIT70wweWIr4cguGe2u+IJkcjX0Sd6Li13EL
bNnAcwdHwJ+mAyNxf2VzFGfmybdfPWe03atzBZYLfQHAnC+ePMKx++dbGUEMjy0tD6KxFU65PP7J
slfMgdwKB7Ki5Ztr4ZmRrUL3Zill6QhqN8QSDU7I45LCJZBFovRPNnOCF4ZxDn/l5PNE7Int2tzr
87McMk+D/Rob85Nf15zbW193H7PemYeJ3P/igss184XPvDHLvkMjfGmLv/cWtK5KpwNrmGHNEMBS
Z5f+tHORpcxsyAOX8rawZFj4RkX9VFTX3QDXBPk90VbrRTj95ICTYKEMaUnk67AIXZU4T1RIXcWH
Ik/q2rzj1sJJhXhgBjSgegTMFwpSaviVzm/LW3pNl7oE7RLzGdcHVY2NYLz7ZLs5/cHkI8K6xmMW
s95HXIPDXxPcpp6vvGEvM2XqfQ2b2/eapXOhioiVY9WBLgggu9LK6U4+/9uxHSokSQtLDTF0OzMi
f4ss5lNEgxwJUAJ+wwUjNzhK5D0Tuds37N/NUq2O3Aib3I7jkPvLcKLMliW40l8SkckoPn185YpK
mtaLUSV/844hVt6KUn999sMLTp4s/QW5QZHulFWnwgsYim6RPRnZT8d0aERB+NHbPkPcFjKMoKCr
yLWWmAlb9NjW6sOfYIlPzKFTfKCs0GN8bjD8FFuuIIwaq4irqC8TEQSKg6+kDqso+dBCGhC26nrY
BRJGQLEoTGO4EFeCIRJtsLKbTqhfuYN+WmhntcdSIsuDli0Z4Te89OqSDkkbGe2JlGlGC+gwAptz
x159P/0s8i6I2bBShIZKs4/yA73PECAporiDRmMjz1EFy2GStg3AOvMzB49UGgCVnMyekEdQBsr0
b5coUHMYw9O5Whq2iW4f2rY9Y9XS/Gh5atNiqRLBWBcZvk+dRp1ZFvTO/vfyF3NGHhh/HvAADZFA
E/Q7LFaHEwUGIIcYwneSQXsTc4yEieQ8ztvPcihBqFuSPkH300IcEiGsGc0v1Us2Yr+7ZRM7fFyE
mNLPPthy3t2Z93/vV1X2DwEfAzwquA7WkrCpvcigJBEn15QdP2Zb0IwhwVVyHk7fF9SQeCIGdHG1
chF4YQTzCNoRXZXo+nBt2E8slXJXOM+JMdYC5CDiOR0CMYz4YaxDVL/N0wp78cyLH9RHwMvYw9a2
X8+jF2k8DoYlJfhljvhLAFus/ySVB6mMtHUJyhDrVmsjp7VPgF4mYChr45vmlAzik1uFivVlIFFJ
T7TN7NyP5JUJZ1135FWl1cV6aa6/LAEWM8/BHD7KfQ9f3/QsckXpSInyUbg/Ymkd1nlAtZDNyxLr
ldnstnrBApCKRMgQA/rmmFG+fHKnhl2FhGiONRRR9fH97Egv9yAfOUR3afr8RB4+1q089ZBA80O9
cMPnJV/eCyz5S2i8LSvluS4TZapa0D2P2WZmYCNkUsF5aoaNguMzb6+DQTzmw/yqapKRuQw/bXkz
++1BSoTsM1cps3hiNz1qMfCmmloL6G5Tm1Ie07xIadQaIEkYtU2qEzxJCFcxsBQqMnur79xV7Q28
YJuM3ryqvc69SrrlUkERxHWGik2Scrmzn8ePNZSZJVnPPZO2pRZJVzWdkafP8llBRHstxP6o1Ysp
bJkHnmsiHrt2amug5XHqwq51qSsr+0fWWCE2WxKbEg8mXuVdNGuL8YfS5iTL8pDwKnuc2Fw26D1K
NVNVsQw68BKc6GG7+uFv1K8IND8RxUGADTy8Nr09Mo0jWXZGYLXni1zMKsKjnq1G/6FipKFmh4DQ
hM7q0MT9960Fh7REErrxAQtZYA5eVIpIYDXN+LqH++4Ouc0zsSNHX0yrUiHqL5lig+NtLxkZNanE
ttR4mGdNJ4+kGFYPGz1W7injWXH3KYehxHl2ps545xSRp0n2AxP81O4rLH9crC0O5OulbyHi4ZKA
UtgFq/rFkes0XOyvzaX9JTWBSKrFFrmiOp+vbsx9YRGadBj2IKTGFHwt0uKvM7Q6sROc2FwVBrC3
g+bwVrdy9BrspKunnEh6pAl13bucv7R2lZLJwZtIGCBPscDoNVWtw4xRikAxEaSCeu9Ia6nbl5+T
nyA5aWsysxBVrtjc4L1vJRjn5LJ2w0j7LRPXbiGaH3LmRApXMLQWPY9obTqS99NWQA8kidgk58iJ
lHJ87frew7XG++fBC/7GhNpalI7kk9MwNfyMekSuDa2zuWgTku4BgxjfkQT4RH/kpQYs82HBWN/U
RanAaZsc+VVTMI4BOm8jTpQdp/HHONVfxzHGe+OmZzPMmYvlmeENcv4oZu8D33gDw+OTLPoSsH0+
d9chb10asvX9IK8DnEnEgqA8/buJ/WVOAzdBxhH1pmxURzXif2hoENvgk6OVP9K5HKTSU8CxlSO6
f1I2RyaAPQjrt1a2MdIc5B5oSS7QNqNwNWpicFaSSGEv/MPZz/Wkc4G6QmzJjqdUYZ1AkxLTQSQI
/kfW8ky6xMn8nUnYf/OTwPAa3Ou5kyI3G9uyvdw8NOOs0hI2geEcSJlr/WA9pNKmGAV5Jesh43/v
Qh+f5KBA3G1OBttnzE4rEOVZ/gVV7ckopGQilL6I8RMjVxm/IObZsaUt4GV/ajKZA7Y+BTXQDKXl
1I89SvJlwCPR1PDFDNo3WHH124jYeQQHI7qiBsBs0ekKklH6yEc2zsAUejP2kXtMv/bX0wTRz63A
sqBcs8A0nxb4TtUHAplz01Fa8y7AKKpoOTlSIP1J5dnGcXsW5LgrMDxSFUXUDVcF2g0D6aH0BRT3
rlnXlBKJcXj7AiR92H/+eOQgY9tiaWOVA1piHW6alnlTww/T1X9edmctf5tDXwDjJ1bi17H353p0
20D3+1Ke8zXYz1QK3ySMi2U1U8ymIITgvDDap2beZLg60tKn+fsxtOUt/9uvtIUB6IccVrcEs7t3
k8SEQyklmnpHFR+qW96Fymn+YXd2JiIBR6Yr9NzQs6J96Dd7SprdKDYVW9IRNWUweMt/aPX3Vv3W
jYHQvPVx0wcnxV/Org0m9/gliHUKuzET8MKjEOJw3zWHucqfxZQVIyCWHbgL43ljrd89xULE+47x
sPuk86UP02Cztpqw6rdiFtpZHXxATazJfSNmhCp6OhRNiRJG9KAM9A3J+6sSDXWEO4Vkb2pf7nZx
0GudEdsPjfC6IK0vBTJ3PJpFH5sLPKUe1weuhY4r9QcrJHqWpNKNWugVt59/aC8tQCd7bpxJlfBC
NDHFqzG3P29E97wB2M7uxiIKV5FMQv8Y2gnCyBcSPMlHhs+BKzZrIrGa/iWoPg+kF7J4LbCPMT12
9CX2t/XtVa02fd3kslih2OqsWhK0pgBjjURdgKiwrLG/dnTuAJcL0npxfgrdsl6ErYCvUUnxUybb
HcPC2S6onVUiiBYQ77ovje/LNG5mDcY3QUsu2pXJJmXNsDWN67B4BS3LLjwQULOFWS6mknj66JeE
kzjOh14pFIxH2a9hB+qThsMZufDqgg+a2Qc9/aF5IPfHkmUamJWA8+vHHjhzaakz86S8ufvI2Zw2
uNiKZ252KAKPCsnllHmKZpf+8Umc0kc51Xd1IC3M7QymRPi99NNKdLICmmNumgZLTxxuh/5TgyUN
m9ELLAAlfJcLLujuDke54m449C7CQ+GmgcRKAV09/ZdbJroq4tiDHARZzKcxAFD+QJ4mg4hvpBTS
xykwzkUGFNgpVrc78i2nCsGhzu+r3Uo8ma+1bgt0WxeUGAgoZSBUBteNIohI6PIHwIPqVWl4MpZh
9eAU52K/dakhjvRSJOsplQ6oYOx78g70zQd2r7xRViFAIIoSzZki1cyhTJGIloxE9015I+E1mLfK
fR/GwpCh8V8E8zpEcYXxGsy/O2AdXbi8XD9Fj41UlezFzVsVLpIGn481sun+pLy3Nr+I17KnrEQ1
SIV+Dn4Nt64kURy6Zwhi0f5deXMXctAYS4bhNbGzTmIi0DXDZRAxTN4cn+yDpLNthtc15Tbmeym9
CbIWoCFpnZPOMKHG5wvG2SNB7TYlmfWBpoCbpC60CpKxQuw3LO14JRFnsmxPw6QZQ+GevfQ0duP5
MOtFkxG9AETYYell91scLcMK1RMKM8rteh8OwkjkKzMBC2YYssuBLQdvOWDfHn4m6XU4stskRfjt
Xvzfupy9qO6S9q0I7zGElyKrAGOVwPJkVJn6TYUknlfoZ/L3iObPDrP/wdnQod0352Z3xy8rfTbm
HJJL9MQTjegzvhC/yuz+GRpS5vxQwh1xV8nRN61v0U2IEyo2btZVFGWY675VlRiD55jpZktdE6Gn
D7wCDr7LuXhBG85OrQ7HJzfDHwzDyZGMJf0saDptuHZ8Za/vRR+GkSbSdfvUb5EUKf/27OF2IB3s
hZmszzWgRHRzt4QdPGZURRG538Z/3OfgBoafxvm8wOdoPiHdrXL5FTEktYHjSJXYrBSaCo6+77HE
aLvyYmDUPNuRnztWSKMyyQWuj/AYF/GOw/xbDvNPWU6pDXCD7fHvMX66gaUVok+joWjXXS8KIv5Q
fl20I9w6eTlUgP+yKVLl/O5hvs6cEmOT28V5/hYfAEmw5I7R/ZJuittKKz28KV+/DiC2Umztrh8Q
zj6hrKWnR+iDE/Z9cx44EOwpwvX81eNmOt//m4CP7/f7t309CPxozEWXcIhQvRMSz+1SR+Drre7w
FfBuqirKA7sh0tYRrqAUJhOMRGQg1o/SP4dsK3YKclFO++Y92q/VYvSBZhq8LKhEfRfoJh7eKQ+D
Bsz8+Ndq1Xa5JXXwRu/8IrVlz1zJQ+0wGxYlM1YA0n9OorcGoQ+9Zk5HpHmV4Gnadxc+eNZEGbe0
heLvQKu7a14KOoubnEM0UpSawJq1fygWgHsF2fdltYLTxMyibrv7Dxh3l3foclGJrnLij1QmgegH
Wez9jdJpP8V/RB2sQe4oucLrYoAED4SIhzZ4nI5qhoOhkn8PMvtuJ8y6kozYTe9w7vH0LWdfim16
Z0WOc3RxJZAoFBO8q6mzDSdIG6ORJt/6qGQZF9KRa9vW/yoZPer8DkvwyhxdkadJX0ePlT/dMsMi
JAS0zT1cmKDyFgcXmHhhpOWNomtZikTpBCGmVYrir2sDKxor389QxjF9VEYdVSL0Q9DMS9UfU1Gc
UdZJ2x8ciLFzsBPj6BSPvL/5ZpS3zBhOKbAo9ftjVrKewubXjPPioE/T2cQxpePiI5T8OEMbycqC
7XRmxCwG9w+RWB30Q219QTjAX2FoRJouzf+hG4u7OtPsHWhzkQ1sprM9Z4rdIxR1ppKgO10aaf2n
IOi7g4xNMDwvwpq4r/rs4C968JZ4QCsLH/AADsWJmEOdaUhYQWYr0ZCICmXgdO1J2xUBUbl6lKbY
Pt10zH9MwE7Z0Ynp5PQKYaTzFl4sKtQrRlEjHEv+6DDqjlqiXSWZaDZnz9Fu1oyreAwDLoOk9Rfv
N13ihopOuybu2Dzhg47e3goaal16SwIwD3bhKat3+XmFad3sXjVeCogOCB3ybV/Zw65fFNnwfXQO
V2cB/uNEQqvgL3nfwY++UkI3vvwZbHadJLmyQOzZhaCLhInHdsbzJO9Z0Ei+XQ/7b+f9D4Mcwuoq
mcYNBpbzyb3duUcEero6ov2NSxLx6COyXAv5tWQxg8+jIfOI5iZiL9iMhYNIP5HV/s8Ly6dmTMTr
ZPyJTkD/6sOd+ViSM5qd2zTsH/QwRx/sNChGcltrFeir3ppYml4oz8eRLiWP+Hx10syz1S7pbbp7
DJBI5ip4DrgliF0858Xmfy30hPryyPImW7IigqfNLFfqQQeIwASDbSJd0RuOZ4revxgwAUsLPqEE
VgnoK0h3okdXzMbDCFebchFMeKHXdxqYktLdFxfxXdXMfgzcHGZ6t9VvklR0oh4rS/zBS0FsAFVV
9AUd/5uz2N42JhLM1+D4pYn7D2sMtqQ3JpOnK5mbguQS4SoRfa/sIU62MUl0vb4Y5eUnyJ/2ihkb
2ICjdPJdul/H7NoEf8PYM4GPjcpiWRmq8HoGwRhZNGhKfbtTFzd4RTTl456g7p6g6dKtXxyJQ6Oa
qgJEMDhVHbgKIW3awOgC9qgcW8hSVkdbS1w85VScM7qAewYEJ8rDNMOspM3X2dsWDesZMcATet3s
QtbiEyQiQBMhMCEAhzmGor7QhBlvujP1rsBnnvA4O5qG6Sm6nlp6ctfIlA0GV5hQ38sl9hPBOACp
Ob3THwPAOlI0Nk5iYe860dFsbmSA+yib9tgUTzBsA+B+C6Om3m+OMCku2TT0JdX42IgqdX0jkxP0
xK3597mkuPbt43SKTQNgp64/BUzNaCw+GStnWLTyKICT06DOrGYKGV+cWLrD+02H/T5qMt4Fz+A6
RgkqrutqQyKxClJlw/MH13oPXEPNdgt8o2A7myKJg1/qn/7JxwcNxFyFuRXE+Wq9tlMoVrcEx3st
8GzoCCTTjK+9ztERcp/FmpneezQ7gJ2Q6DM+PaWHEzCW7NhMfCcTHWXqx4PXRuRDkhoPE1kMXc+a
ndOzWxrNi1f1Yo1IXFNmvFY4NV3VAb6EgymccJGr+P/MSDKY3sqfhtc4/ALxpnOT5XvAAZupiCt4
ld+tYGzoMqJkVL4yv0teXT2ivMRrw004AfyKWfn7bhg5kvmVTVP9lBAT/YIkpHf9kPJx7Xk1+dXG
1AGXYHxIOSqnltpRJAFtXFKq79cScVRKgKBVoz9Te7VQTTbIDdSUtQ/FXbVX8erkkQCEUloUKVD8
Tnr2w3AivLNLKTRQK+bCP10ErypeThgkdAL3Em8fpnd1EuJDG+xN0W8JckO9sJo2Kvm/HvGrG1aX
zpVMGh194rSxdy28KFYAPSsFjh6cnUB9w63ZCJsrFNTjW1KkI/rGko/mD4DaQUD856Vc/4QOkDX1
k0X8z5vQvsLMgduFzeMwNOQiw3OMUFYpCHB2H7oYXOGTMeKpf+jlyuc6ToObAhuUeYYlJLzzseS9
iPGGh5QLW4Zj8x9rKWPO8zWe22UM4qwwIEO+jqJfszqowNy2FunoDmg+rkOR98MeT8idaYzdl2xu
ueOoX/Wnec8A7H72dws0Vd5IOep9MZlx+j8NBPgdpModJba2Wf8R82QNsnLCw48NoqIu2yoSQ49K
evRsHaZwbzgQoHsDrMfKoJzxPEg9RdnlQS+EuxtAID+wfjToZHh4i4G09v6EeRwDqtSSTnidB3X3
gXTX8AUGTxPNd1VJl8UKibqi75cQeKAuKST+c9c3J5cZA6zZoSQKMuGo4R4GdxA5tIL86hLqlt7B
5RnsqgrVSCzoecXhh2otbUQ3bBoB/9rL1s49SJcxrEs7zTcPcdBFuRG/im5ccNmFjSYdb8x6SWNC
k+swcUsJizAB+uuUxmP3f/1inzy3FGIqIzaRJTJzt9GahVhrGbCmLxjg2jdcLzZYLmwo99v+M15W
XvUfWzlX6t5d5+3ByPuX+DEh/cnKhfbkp+60UvWBdr+VbpIe5b4TZl4XYcTqw6iQLIPpmd4xr9hh
/3Nr874IMai1Y2VtFcRee7TU/m35q01Wx1jz+jqVCnA5z7kNvUKJwg6o8mdE62+ONTxRj/U1M72g
ko3qtcj0svx+i8Sxh7WSm2ljbQ4/ZBhF4Er00dWRGc8REPQwoa2feWaf8O5eTJduF1i1dK9i1J8K
hOOwCf06t+Xkxk1mNsPmWA4s0WIco+44EchhYyYo2ssG3IUXC5MvIDlqM+WwsjxGr7HEQtZXvNTB
qtbRqTeJcbed6jFuwfIcLnV/Fe9yzZf5SA3Ti3vzTT9wSKaxi4KOcmrWJHGRZpo47iCP0cRFue+F
NZcUzJj3xK2R3LClATSlwPC0mgDXosA3wbz+gPgatSujIffzJ3JiFVA2iiKt32wr4Rc9yQUVvowN
nup2EYKa1Aqi+k+GUBsrYQzMO2+dFev2rAvX+bztZspkONf1A920ljba/hbRmtBr2Y4yo+qFj3kg
YfD+PtHJmSfIiFSe7cHd9kyziKWoc5bBL2JS7YWm9Zxc+QWESJJWWYJtrKWVFaCmMLISD7thip+g
n5F59gIufECftMxTEgcJbVcrW0y3tYTuMIZ+xBaTTM0mTmSdtJhYBoOOuCkZL1peL0tuMCAO1JjB
BcGb0Xu0+k2dKDgk2zOiV5wZTbOAMYBy/8gZnPXBqRoxsxmq+8e1gmVLMJkQjALYcy0bxMKwQ8o0
cergULaf+d8cALwbZSOEwzr/h809X49CnaDIOMLQt2txxjvWF95nEA30QA9zRcwYhBqwd32E8Yqp
+UVZrYbXpYA6EjGtBQar3cy+GZJ/unn+qK495cFuKpXiv2b0gPuPMy7glTVhipCTKhlwUV1znsgH
KPL8cgt4ervYIJySp4ws2YHFk31SQwbpWlXzvzuuzPnd8BfFQpVSd4TClZm59GdoBUZo+5TCNdPE
u50v59HcI0fzk8GanRZcZbIOqTa1LHE1JmOFEQO4mgykpICYoIINL5JzHvR2Ssy8JKgG4aWMuZif
KBqHZPCz24VIU1SneQ2j4e3ujN4Nuu8z3+UEWvN/KoNSEPXCPQijkxmJHh40sLlZ1JzoRqy0gGjj
pWqz7TAk6by9qOPFcVsQRldpSD1xqWWc7papSsbHY4gm0YvBVy1P0X3PnfppKzqAwdfgV7icvp0B
6J13NVfxzqx8JhYTIGb43Ph57uGeu8kgvIneohQu8g1rQRwv5x4ihQgJWMLj5QadQONWFp3FP+ZV
351C921uylfUB+8tiYSETxIauwTDWtWypOubm+dt07gkOnCKhiPAmHR70VtCLh4zsYpaHQFUwtxL
oBJ8W6fIPl8Cmy+dulwlsZ56MOT9dQKBgjRFStmtZzoMLAC1f/86r9X9zcuGvIEgiS0q8rrRAnzG
+uzcD9B9wQ8yqQ9VQjPwwG6+mMmgs6kRfEX9wNJcc9sxexAfQBTuDY/G0HSgbuKPOm8aM4XgUimZ
JHIlEDUk5wOyllLcHiAiPWc1y7lsxFp/Hs+rHP8kvwSyO/Zbg+tnBDBAych04upcYgKWVc4ZPqw2
sWKsgaoZz2RJ/14px/AsfU4ZKCOdgbvahhJPX1H/KcTXjRfNN/MgsHYPzHAZlGknnvl2TYVPTLK0
4pjRl+dNb2Jbm8mueefv6naDIMZw+Ulun1qjgNd9mOf2OmyCX0ktkh/w57HFN1kkJrOCZn4oyHxE
EpQj0kW6VhN7HV9tOjb8n+s7farhytvyIyzz76aHzqDHroMcgY4gHEYf+eHMyQAe2jinA+ad0MGB
z4ujcC6sGE7XM5JDgR0UdSY7mawSDHD0FWQkCEWGL/jE9cghke5q11Puz6mhMEv53yG5FZMX3TVv
+pc4ZoMhVDziM5RqpXozH0mFXwl1TFfETT4iEzbNDbZYH9A2ZyqnLJcb1S/5o3jGmUQmVPsi87VJ
Sf0rRm7QMHAkNeiVpB5gIkfqNta5Zj1RsvQ0emxvAKEo5vwXWie7MZpHx/P1CKZKwWL6WbPXZpW9
PjydaxuQKyKerPQPh74fvJK2kR8av/yfs8jlKTszCUIko+QmCGTmPsNE24uFVX7bcyBaDpevBKOo
GM6LWNOcJPbvotLRjE96FL9JTgvu+B2uiGsyW9A8/P0MAoMzCka9jAHik9uI2T0OrbRpgog6nN0y
YFq4lxkjroa3DEWShO92ZhVIZbaVQlzZ/wiZv6qt2oBuc3uUieDu3DFrCpQa6JATTJ5s/1OKs0qA
EPb1e/BghXs6ilCk9E8norAFDgxKlcCXbsSXH0Ob3Tx4AblSUI+drwL5B62h15PhEqpg2JagquIJ
TUmtvWNTc28MhQzwm05G/VI8pzxIpPRLJqzXE9qgPirKx5zxF7L0Bk2CA1df5HeIlH9yIPLwSdj5
akbKBS7DKiCPbJDsguoxp2929wbqi4kwZf2h6/P3Fp8Zy52RukAO/zNSYXCQC7s19IoNpv6NAZcW
ZnXuWBYhlIyfjz9vHWh2H6qcw3Lj2Ak01yw2C6ci/IF+zQHwVvyeNvbAo2PieQWGyom0Ano606Fr
C9o8mSXga4R0InU2V2XynkOkPcuFQm5KRVdzbtZ6Tu9ZVev2DIE8Q3azNvm3Pp9vn8gm78FtRNCD
cMr5NGLRhZ73SxP6bssSvIFtRoPY2slowd7UA5IbKbPp/UQyx4CgDWd5DurbZBcJ+hdeBTomuL/6
p5wHjgy81tvnfbz6Pn+pMwbGmHiXJrmFUHrSYNWYUffkWrHP1u2GwG839EsZP1UiD0LmYNoDaegn
6g/K/3k1HxNhXndCcApibak7AaUrCM7MzaSUCPimTJ4rSEo828ckrP6ploNGjsjQy0NKa8P/CasP
DmPief1m7x6f3IFexKmm6XQz1Fxl+/kFbZVcT6tx8dUdLNsnzNwV9WFWRRCDt90HoskmDGZEClW6
Siajbcrm6W/MVrxqx5kq1ZEJGW2p3+doUIdiCVS/sWLUq/Hd+iO1aAs33dGbsvHK1cYLTsITeF8U
q+yhGRyGw6ZdZxtj+1yHcGLZMrev0moyd6YbZLqG0fejPdS7dKvikf+9b68kk/wfqrJxiVC1Iy/A
x1IzU+fkVlbZAlljBcVbo5e1PIZ64B8QSGXzOMmN9002KhjOnzNFEb5bWm692Vp0gDc7aG2KLva0
zMmEulk11zvz1JNMDSshjF9R1YGJhjmfPWA3YS0LH3QeMRx3nVb8Cm3r28guqP3+HPU7FLWTl4No
IONIsgQpSiKd7gN6B9vQxVh3/jNRMlpRGFfOyN1PtnCUF52g6BLUKtDtBwRWKVwLAl7CbMhTKnMw
x8nvFpIZXjt+MVx6uCoL/f3qNKG7+oZjVa3JEK6xOT2wohtdKZETiiCoS/JMK7U9/aesl0ANyoe+
tTvGciDfqhddDj44GcpDbS7E1QE1BA5sdRNTRhp96mvvCqsrZ+GUN9k8qfWXzAYwAeOvgtWzUntJ
son6xsE8UkW24HVYEZkr9w6vSI31vIaCy/h6OLpT3xyB0IPLL3yHs4N2ZtF23gZ+kbdnjBjmjnQS
nN3U5XwIDYSxE7xB+9C/t+0rbG2X9tNv05dgWvy1EJ+kKHbJGDyMtKyO5PJYUAjydlqEQWohJVKe
7WDFjru6MSawjyzx/ZQMxw1LmiO789XSIs3k2N4zlPBA7LVWjtDygSpSJE7EKkJIaUlGyPDt5RrP
RVHfNjDhWQSUiTKqjoCmn+zixFlUk2Xm8UsWijni1HHYhEIDrg2jjzSisTtHY2UKP5e2aeGdcyeT
rmEZRUeFYabOkLC+20N48ja2VRkkVxAn2oO4yzkWimiIj3whaMCeiPvaTqnabl20lh0ea6aaljUM
RQjw4pxgzeuZWAmE4bK+dt4RqJZ4/OAvUxUlImQajdd5/i8H8EyA8wnX54k15xDSOkkNJJLDDtnB
y+vJe9tHkPYsbfjUCb3+1D819mDdA70QQZCR/9l/Je9UAe83TsYQmvvOlQjD8ESedh/f0YKW/xHH
ytqRIs6ZETaDjWlm9M2fYMw9YC+G1OwUovDjjpQx0qv0LBvTc3I/9DDHrgVaBRLbDzdxKj0dFZYH
7YePW75nxtgFJklMPCEDlR4AJeY5qnOH2pG3g6ILX9ehg35PxDrGDPIuB74qN4JPQHaX7aeQ2XPd
cD0jn3OXtqqHh/gZsoWShRZNwAwiC24xh5hM15MuUyaGfawSxZwqzc4cGgWVd8Ep0VElN+mCNN8V
GRsg37cMXtetE/bEmXmbgjlSJe9kNQeY7KRKA5y86kNOfrWOuSroCnVV2efzlW+8/3bN7RfFlNpK
9jVUs9HH1jymZonMnx+YJ33qdwcQUQ654J4AUyH+ucdJ2mxwwFyT+d5C/FVDpwWESPoogTDyhUux
sK8DbWwjUfRq3yTxo+eCWXt8umVtrXHBHU21p4134hfM9SL8Iw0gAYzUb94AUdyr5NTshOO97sZm
h3XtmtVEcDDg7Xakd+9ts0Ref5bn4UiwAuM2/NRGp1aLFEbqkcb5Rw6X8EhIcVUObbj9rXVTq8ty
Q6ou3mzo++AEHIs65Kum4DQxf7PeIXlRqY85wY9J4WKwM09BI/qbG/bqJp4bsnU/mg2j8V5Tzq35
j0XpDYl+QiAdAk8/Z4MiygCA0EFSd+jWwNfivOpNgbPJ9MayKaXpfLHzifsoFFSGx2nuG/oYX4ul
k4xYBmW1EbQAmy+gKl0fdqV28zJCqn60T9nqLO+/nYAgf2vj2Hm86xa6BvJMMk06KMcJROWLHqRp
IJWc2xlRb5bN/eGpBjbH+U114A/n6/1QHycNej//+yUtP2uv2Ru3OBByW33aopIkozMZTtfliy9m
ch8T0ZfQA+KNciYwkH5vBr9HOI989uguZc0nSM/7GS/f0iucn69JRtCmWiJwrHbdPwg+zvHvIRL3
t5/DEqp4w15v8lQ0Owd5QhMkjfT8EDRGvxIIzWO1QJ8+mcTT70XdZ3KH/tfigqgbNsetx4MhiuWu
Hd6qHkqdpIuIRBGHvmd5U4LK97r+ehnVrBo1N8AdrcZL6VvrhznNgX10YrzrfEA+HhnwgpmVII7z
3nHI0X5dFARCnjReUE54fJdrfG2cKKH6UgZ1ZjPN3NYgYNfSny2UjYlHPuO3gAaHDJi/wkDHFiy4
rXzz91eNCTIbP/T+7PgByy5Idv7034h8ZD+TqiDgI2GB4JrbS6ng2spmv20OQ+tYDevs+hUon1bo
SkWucHO3M2TMNUSGatOjx9SUMw2zC30f43LyXJ6Owoz1phKJtD548jw3EUZnq8LjaG8YR0IbUVIr
iNZK7ACBMdCNSILmTZLV8yASDTu4x/+ajU4HvFH7W0fWguVY25htHDZUe1nOh4SluAnh7gZYsIsi
6cupH5MrZhvZweqBI/hYMazjNf0HBto9767jqIGtwbUiJDEXQnseeb3LAqUuUBRv8KrZ62u061rp
Rg7hwOL5MWKw9T+mYw1VN2xyJ8v53pD3Mq51YxIBa0VKbTZH5yreinEro6Va0e1Ru4Zr9t+8Bgt0
+q4mO7ea93otNn4ULLjC2MeOnF2LFqthXa2lb3UeNInhXYgnQZk4r5nwiHx73/WOseYZU+BLVnIL
b4ueuW3nKAoTPYWoMOU8+gOyhQ1f9MrqflBq3q+rq0HFpAlnHvXUBHFGru5gPyUpzbMPYTENfJIZ
5gNH+Mu3a0lGpfhyncJYDbwaXWa1+FAWkq8RkQcf0V5AVaENM2cqnd0tFnzZJltlmh2Buub45Q83
DrcUJ9OBvxQ/IZ+WHWFEStMFmSn2WdRDDmuDB0S+SkETZ0D3Snn2If9iDfoKpTIKms8xu0i6aIQ7
RJMQ+reiEQMixTUNgJ1vl8X+eEdaKi15wM8/MARoorWiIs6n37hyZDwgxssSmo3CJoBmLlVG8+sv
Yb95RpM9dgroCOIOrFI5RFKaGkUAseDvm/t0ZF/sBk54wlQMg9QmKu+oeb2koKNFRr4qrXDhr6j+
xU2qcQ58TLPJmdl6KJztS+U+2LlzpSY6bOeR6iSDDVkD5mHeyeBOmWLh69vOdm5OeRjJD4sR8kee
2Rcxwk+0zKdfQf8Cba5grnQlh8h6CNFmBSaao4uDIaUCXZv+9FQhcxAqQjGzeFTlP5+wo1G1AMFe
1uUoS8rEMb99RUhv5/nsZNDl61BPfH5xAYEFRvHCyt5ddqUPvWfM8/ZXLAgRV71Gt8HnwZGLQHJg
ejQ7Ac4eI4327c6FAFJ+PAWodvNeJ0JWXi3pbLCwOKrwWPhs0XpEAZm+kzfd3nt2oBJBJzOgMUAm
+ukzMgqwOGv9UM0Y10B60fhwiS0WAG9Xj8YUgKPjvqnUyoJf1fp1qAP2ShbvYoj1Ok20byteSZKV
6OkPpoRtQ4w3S5WWOhPyp0byOyim+OnIiEunek+V0O0jpJKtPZSgMi+sxsIzs0VE5ZF1Rs+M3p2e
Ca026/1ABvwoRmH3gBjS8zwO2kWiePAPUiYVdyoH9jYX8AtPKqceQps8uDiDVDmhWPwR1DbS/l1Q
+lIA1k7g/LJqMu2TDYgN5O0vAu6+CYQgHph0uMYvlVvrxhTtBmyL1SzYDvf73TB8penZLQgjXS/6
Rw/4v7WWBeXQsJMR4JyKSo+ILGWIw0DZwhayd6MOFP4UcI5zLt8IrwO6ycAkC8JkcYcLggQMKOSC
vefipJQreNCFcXhJ5GkzHcr15jtLiUoIx9NdxTWcRZV64HO1SImXiHPzn8unehS9j3z8IAONWZNn
fsyppi+faw6lkGZ2/FTP/xIBI1qBZPjva2/4WfXrF/fjRzsfwOox/Hb+YiaXbZOgwQ40MOle//9S
xSYu2s0iTrkQ7QjKU24ZPJfCC87VPrEkkeg2A63JFt0ZAUkmETHWehid9Vt3gP3f4p8e9kb5H94Q
oDKGxC0oC3Aj25/YVe0+Ze1bw05xl1FFTicxLdfvITGjoN1i8UjWdJHZFh7l/XMgEwVVvDPGvdmT
rDVkAtb9gOdxdHd/GusesTASkraOkFzuD7MTpngjZgKe6FH8KmJXCFf/ZQLAuq3otP8SPrwGYD7B
JlXoGOsB1qm79dlycHCJT1QDPFNOB4aIIifIFyYj/bd9F+TumZqhBbYnZHpgbV3cdfrIDu9s5Nas
QVy4ZhZ1EK8t5ZVbAC4ju4FOdc8kVIxo1sfoLP7gw5+HbH+/oZnmH8IgcSO3b3uo8WubtaVCXpmC
1wKULdIC1zyKzZeUYZz77xZK4c0+JcwWy3v5tAqjbqJRN/sI7hOD49nJQw8DE9FrWhIGbwR/0IOA
c5wEUpPw0hLpdV6ZR0ZSFhYJbOuNwkLOQ9tnAY7CTND3jtdJWpIEYWe5jkKOvQueVxm4pWXCz+3j
5cJ/TzYCOPcfveA/+1yukAD8GkMFvBsVgjCEBK4/0Qszcu9kFJSumudb8P6nC60IXx9UL0HYUZiT
ROa6m3jOwUVMVYBcYZLSTsnxpWtymJmQrqMsEsBCmSaRzJx9zIZ4nvtUL4Ni2OSgeYuMh0xmB+ed
oy5NVnfSdSmAcJ9znDW76gWck5+NgeyS5IS4MVeg8Uz82LboO729YB06r8jpGk32EVx4/c5pKze8
jI39dPgUxzv3ZUtQAF6QpWok+XSbe0vrXPGtnKXTC7Y2lkiXDL1WGCrQGgnUaytWCOzs/8qxgyrz
K5A26uIWZLknucMJk7UPE1r/9uv4Lmq+Nl+Jo5ugVeMvsPGmSMT4OHCHcL/x98+ZMojEAj07fW3l
oODl73NIzVP5iBiGNqlF9joALBX3YwTQFQHVzmEBql+07CAa8kWUWc6XjPHbjxqiLBjuQ6VTUq8j
ljIUTZBTAJUc3Fq+IDZTFXOa3JKdtQzb7i+j4lRBSMx8/kMI0p1vnnhA2uFEkpICYQ3P1tiFB9HF
qH1qQgCLZcRnAjsySjLACHiNm4ZpXuDhYSZEbeg9FCqEbBlt2aAOCMheb0Kg15DsElG/goUG+bcz
LR56CiMPbr6wqXiREZM+iDKXoygG91T/SdhqZ1sUWutx+TePfH2cwkQu13MH9At70uGjOaySpPGL
8qd8E6/QbdIxyufLyBnyOIT4Jc5ZXOzCe7VswaIsOwQQhvC9P8r0sAIbRNmb87BLVz82VUgo7H0f
650GdM9pSjcKWbHggGbN6CR1RcDSMzBV5nFr57rl+/Qc3DQiczsAE84PkaEs3qXJEhEV19Ds1zKi
skGi36yNEmQOynccmb8Cv/7Q5VXxA8gB4hGcHKaMACQRFixbe3znhnvVZgfCOhx81Q6Ai5p7EqdR
qGXK2Fq7uBF/leLHEpSif2ynytW3Q2dDCO08MhTVtan+d+H+dglc2xjyaws7C21eOd6MVDO5XiZJ
9yS1VCCi6zPoKkKJYvLKkEb/Dt7wKOTs1LoLA3qB14KoWNYfCERqNzyHRawY9sCiLifIqLf3xFFz
J1FL+PXN8JVDAKaNTnpVvf/XZqNKyfSUFPbgRzjITBSKrKG3aCa+f0ohqIhrGSpW/zWVCCpHdcBK
LdOwwQbrWPkSjZNSmU4b09FptJUZaV33DW0PbhlhhV/hA/pj2BJYtDf3KDG9Qny6V9ogwzkDiStb
QAI1glaV7+jWl3nDiYs/X0PE23jwiFUouv1VlOac5jk5r7qxQHRViqoGY+S0yz2A8rK4gELMc2hv
2s0mUqmGo1+HEFnfQtmnOkFDIicNQyh4/w0C/HsjFmbXJh4KNEZKpeK3+GJSNaincXupyYQKIZny
tdXNX0L9TR8cCxJMihE3kJMztKgHn3elf9LNhRu38/AjNBEAVDlvEn+9Nc/bTEkke1gi5xRZmmyu
/hMzfvay/fo9rBgrAvr287Xbk2o8IhldlAvY+sn6eFjbSTZGBuWqOjj/91sSEjJ6B5+YOsZDo6Pe
614rLir/8KHReECSNHq7czp/P7PLJFA4C2SbaIAcurquX7/MZu+mmkad3ZT4gVAtNpFNikLsysPz
82fh4cpwBuplZKxIyCvJxKlZ2x9FSMdh/HXTuYvqjAqhQeitZWkPjN8d2X0Ip5W2WbgC0jRBZXmL
6XR5smtPCEMGnGl8BbY+ln6LtymTJ9W6G3NlZ1UtVAKm3mG1FWlLtd0UVD7RMuHNStravEzDjN9+
cJ+jga7OrFn5SgPn5qQ4CZwys70st7pzYXRUtBExRGNHbu6R0a7uei4eU2/hz6EWwvpdY+SymPop
MjdUYoGEWSRyJxisvy9p9WZHyco05a1swMI9XNI5aoj8pYXDHF4BTC3pZm8vju1xf1G1sE38Q5xM
SJvGCD2+Q6BE4u5ufZxZ5ZGrTOms0H63mOJUBkyojssVya+jNeMSwmZQ68J41WH9vwLb4JrGwR+B
Kj8tBZh6cREecWCkl53DlSamXdDBmcscwpBji7d0dKCmXOoGAo6wbD75H4q5rLq5ha4K2TTvrNxW
M2CcXJT9k1SOIuYsG8T9sZerKd0/O71xamOtw1KnQR49LsBYZlHJuDVmMoMQftdi/QoIRejhlgCa
KTY3WRICwuZnGgyx3v7i9zb6cGSlrr9GQTT0vKSjFLk4H2cnSfdPjQbGiF8P5pLIgfh1fcuSIa9M
F6VN0pz1jv+Ha0583Q7IokVe4ZDIc+yd5nHI5fsQwVYcV4LhGG4QQl8dW4kbwp4CK4RkvXMc1qxk
J7MT5qenICblf2f4+cYGpI7qCyYAZOXX8gbsQuACIEDSv1d4qXiz+Ikkp0cdMTX6v19wZgy83JUW
EbvX7wfSpbtn920sjbatpeYLUTVOhXRGavzdB6tLpwE4np9WK0TbgjjzaY18BeoKUbuB9LuT3YZH
yJZPTSUwcTjiaGjV6GFq/6W8/FeJMV90fVQBIhVS3tmi6gy75RqzkOx3UAUFrb2o3MCYLItPb5jT
CFsXXtSAXiJhcYn88MD3XWL99/xcUvFKPi+u/g//ctJChn0/BlYV6pLW8hfcTBjFCGN5ZxqBkJz9
WNZ24sGoVqMZ6k8a5vSBha1aRil7C9RofyobJ1n6Yw05wDO01fKcDnjgDaGZSWZKFfP3Yt5mQKyi
oLLHvwoOQIO1GgvuauCVaGD1PuG/IYKTwjnUxXAJXqlKceflwrLJynaIqaoHj4K4iHwJr+q2lAtf
vMHC0pM5CTf3hEfShLwCcusbA7OkTdK7TvFgC2F+8jqyzM70YjzVh23z0eSiN6AAAlJjUk33jZnu
10wBpKL1GSCynhvbA9nhFI40Mhil6H0A0eu9NwGPP9ST5rJgHjITHPNG46mk1Am5KX/tX0AlwGKS
6g0jhc0hPtM8n7oPcTsQJZFZqDsi4heiSKQoxMOAkZlLuS9Ix1MT9mGzMWRDaoRENCPV+rcSZU64
5v4AC34+4yI3buNwLVRuiUnsFYI32i7wWOWTksjuOBici5A21WXonyiUpBrYkFCTyHosLdDN4Yzi
4Igq928OhAWQqRPSL769bSzkHwahuH623RfK6QXK8ud1/Lszd+731QCD1Z+GlLNJ9el8BC3Y5AMJ
vTSrAtxI+Ai0v1E3LwUgP03FnMI91bSijIY0Oj2/0szCZV8LBtp8Yz6gi4uzV7hUKWhveXLEuctZ
0iE+lMqyAew2NhlVXYRaUGt0me9HGb+SUCIOZwJYSy7ActO80vUHbFpvD5urHua+GqzeGdJ3DuFY
3X/jXgunRGddrhasJo+rvh0Dc5kZMs3zJiC3A+x1lXEt5w+zCzblc4aJ6g8MgoQm+DJFoDGD2Q3w
hcGvk3f5Hr716B61aBPZ01D4j9Q0cKefOQxg3TVRs4gpuhxKZZnqm/ZlTP/WmxHKep+AU2S/6lGx
DgyxNIUNELqPuYTcsF8m0XEw/HCXWJ6yhNOtl4ou5B6E5u2zKov7LuhGxooBchXzzG7Mgc/235h6
e9Tb9CywlEn+ZMsFJfo0G/OnCWsD3AVpqKrEeHDVf5QbKZOZ+Z/Wvn2ANZYicXnNetOODRPV5bGc
MkyrrMc5U4kWmTtTuGFj6q83YynHeheykNl5HThEzYdkLhnOxc6nYExxp5CuYr7ODt+KYpAFoe8H
bAC0YX91mrXggqtzY1Gv59DHhL5RRtXICLb6vywfwpBX9hTZrd4qCI6CDzHhwKqZ3kZMn36w5gXd
KWHffJneXiSk/w9bznx/IyL/vtKggNXF5jq6V+HvLFARW7ZlGt9z4lTvjI1QV/nerplYXJeo8HAS
g0Nko5EgTqHN8glPJfDQW0qGuAtItlKoSCuVFXRU5EWq50mReELfDmoPkHazTH3Ov5xhdjeP1b54
jgEO88Mbb4XvmJg0SIcvAfXN6QvNvvZZIXm/QMi6bN6SQxfyJOFOzam0DwVg7H8fLs4fbDN9knwJ
WJVRCP/hqlEQm7uUtWMuN0TjPdcoZODrpUvdfDwvjT/VUXP6VeuO03KfVUyUyidsN4qsik8kbjH9
6lKclLHa/GBlDTbRTdUMh0q5u5S7FPtj3qXODgOLjVNNtexaW18JrO47KHNMKnPSIdhtvC9cK5A3
iRkp481jgLy7pgSwWwVWgeJNwy8Olz95Krm85rbwPx/hHPQL4xo5Xkc1T56DpBTLvzGYpHIZ/Cro
aM+8Wy8LZgigBUst8RRBu/TKNnutPnvbPC09hwTgUeYKPTXwSZlaPS3TwptWfXiDCpvNQxNtwalc
zjpCRnecuCNhDiU/JkgeHyj2pwk5fd/D7grS3d9pk6pfJCJmRMIcjnNLpzU1Enq0PUeroxGsuits
12/jIR8hiDLhu1msTsLzFoyM1oCwc9i/VQZFAJO1WpXMUaW4SHJlVls+PpLcF7sg6CQWZPrM9VMT
qx++fq1H1mjgSOqIjzyyKSksMzeMW++D/Kc5RGVi7NF3rKLTKePlMmg4eViya6duih/5lOCV4MOP
ghjvYE9zwESIQMsFC1ojQ28PX1sUlc3UyMSBJ5dGg4vqWsLPXgbMOZiTUHeD2zU3HLB3kTswCTKJ
nxNFuE6zyzdG19828ReAIrA1xrTMYG0puAc5blMOXLdv//4FQuY00AI9Ihx0Nj4ArwFJtxLZaArc
oi7U1OWPUpEhuP1Xgvt3CutmhGxfNsxXIg64isMS6HoAaBSdm662htzQXJMvbcrS2blQmlbzdPXI
ylfBNNeKpMJ8Kmit1hhOsDgsarsgqyrDAi1L8RJb+f/0Ndx5ULNAL45uzWklH5yjE6JYCfSnxlBO
LVQZs8ukHDR05pXpbN5s4zJO4Zffzm7KIrfRDyMEe+lixLQvzgECqcEVe/mt0L7nYp7op/PzEpa7
JA1ZYCx84bPZQUKHw6jeRVuhWpX85uGTxQcQiHLGZ53Yh58FKmFhi/z2+hMZYRrqud0rA2sSnfyq
V7dNFZHmD9pCWmEJ4Qpj5xAqn5iUnjCUMTBUqwf9vlZtr1+z7L7Q/FRy9Ks1cv1jwpVxU/hn+jjN
KnXRlNw4Q1B2DPnxF69eebhDZFP7jokifQaBTERHSDfsa2wdD7Kr77MRVo+TmmfzTv3fFjTpvvvk
JTf9R9HHZ84k72NbmxWUN1lVCL7MKs2CPxRHIOYzsUfSQEr6CQAD3YTh0kK6IFHstGcGfvaPD+tI
Q6Q45nMfejuVplNp0P9w1yPvIUGDTfeAhURrQG3799ALmIxw1GP387S1xuuMCMB4crM/NZPEnry8
D/WOQUCWfBKJwcx+yN2rYRM4kN+OZhEG4P6TW/z14faUYgfJJJf2cjAobk6xb7fGgnwFMcjFH3kh
meElS14LJ287zSeXf6ti/CMSHwrLUfXMgYrLFs0wQXrGX8DrBRC1RLmVj2W5jaiTfOxOjU0S46Pe
jq0LEpv6zZXbeY0JCuTDNPfPedEmLvCgEw8PKIaQpFX/oGAPaRnm/bYhjiADArVMlgZliAAaIT0l
SwkH5AWW3L4skTXkaIi+le0SzZAf3blv5RQgoTVlduVRlluWMLjGY6IHBRKBN+ChZquIW/MhYKYc
aTwebMWgh12HZAVP17wDa/E/iZw4GA2yUfYsOZ76j8f+M+9LVEP3Lc5UGe77TZGPUBeHegJXEaKG
wSr9jL63xxKqHHF0aC4S02b2bcXfED1vLYCScA14Avn7hsNaI6Syu+ZOgnBBC6dUsLYU5GbgpoMO
JEYiBvG2MTaIvRqxZUuSMOuuGsBDkoeZSvgjcXDNJXOZffFiFcZIv208nRuVnyYz+uba6RltsyDG
4PqDseLXCvw+k61HerUU4xAkN8EDR7Xwj1WSjaSNPvFt9D8GuvmhkFAO9YUj/RWRwcxw8rTRuRRz
EM8hfi78EYmMjL7LjYCGPl3TO0yMvgt5XrAai+gIg20zoLMwg/0cVx5r6hjaBdI2uAIiNILiZALl
BMbI3T6PJrchRQ9mCgsvYHrAM3hONkPefvv3hcj75EeZcLMG43/Svul1eb5RzXXZyEnytUVczn+b
NMOy0mIfmnnscIQOUHhMdZWvm6b0VXTjKml+K8uPjNHCBpKw52VPl4XmVl/Mp6Jc2YWW+7ZOIvRx
zASAfzYTQiLjiW3OoDHG1/rrzVLFvvOtwy7MQrkJHXJkiATv2tFuxbbsh6v2nc1HWMiB0cbYfwGo
0WIdQumDYrCFwXKFDcqoNnON5S+hX1tVcdvG1qjifSYwVqcsD89WoVahfYi+eQKhLJv4etvooY2e
yx6UrGD6TF0O8lX4dpCOMprB43dJjwmWeySE3Hu8Iw31HGlaLkZ2vl6f070tclwLdlaTaLLuZ8Up
y3F/zpDF/LULJTCyRjYbWeHLPx9N2ZLx71DR5GlcWq4VbRpdZYIIW97vPwj2Vom6HxkmxnLooDNa
cDehMCbOd3Cb8CTm160OXv9C9WIk0bNW3f+4Ki33W0hEb64Y4dnSy3OyeBwr6qEuPjm8PuImG75f
jaApiO48xBrx2Aw+urCuzLzFbdoHXDGYI3SdV8fOuyBAy4WwQ518pwVZQ4F16/Y7P2k9VizvNb/u
BpeMLGtmTc+q5JoVkqGztMKiH5kt377/jHWCa4i24DY2hMSvXNNxUFqul2kjR9C+xd8Z6HB+gzTF
bengw/ZXMrXdfXKNV59KDhCmQxNjHr4sF9G3XWCkryymI+suzt29nd7TWyMr+gS4Lw2V40xGYn85
0dHMcIqfY48gHPKyhsG7XEkPltmSYjqIQAftu4eTX52KXItR59Pfu87EYwnkDjB56I/XkTPdHoCe
tvV3j+Sd4FTSLJQYagxKo3BTfy1ZKYiKzK8ZrQJuT3eXaLEezT6Do91uQFpcUWHhhtWQv9IscjLy
UhQ7/juVLSF/7r5pTh15Z7w9OQjnSZpZjhIa0b7FLDBMB3HRqTVCSql+66tWLf/C9nem8rDj077I
4WfzHO3E67obwfQt0Vl7D2ylLQPe92EN5GwPndVM1JO+RQVEu7il88uBuf0a+DtQFbHu4R/4fDmF
aZnxb2H3WVABef8j4f4tcetVULSxOAwrvLmv/D+5PdvrRU0non8x6idVzU3srxJJii/hvkXSxkUH
pMYKugqZmcw8FCuiMw6dIRnIGE6k4dgACjJDfpA8nLY+awWM1+SggXD+2gZ1WsQ/u/Ns2sOUnui8
3OsLoZq6qYxmio6RdUb43qkYbFhvrVKZJgpawLJPJBJzGSPus0iXIm8RJYq/2T8N2d8k1dYfHnf6
HRv3R+PpTVJ/Fv16gIGp7fX2Kg78DdQBzJaKi4KbSICcdBs3KFXo0lRi1rNOyWOMZAEyzTlc7bCw
46PnT5pfC0R6dK27cvnIBlw0NQLZ5avEtK3/LEkrMcoQPshCy6vowDqtgS2DKrLkgHHRQvtkZinh
zeG+Pt9k5xmzax1dUSRR5wCX61pKyjf9WRbSugHXP09kyzVLK71UVlS7HApOyui6lj0TK42aWkwl
tY4r14tBSn7ZtGZ9VHh6S++d7EcJ4ACDuPxIS5u8NFWsDyYBrd2miDhqTEsP3Xia3wvwM0ujav5Z
jYQd1VRVcIGA+xVHhccjp5IL6MU3C6QHZ4SWS+qh44v8DkmR81v5CopIKoKui3wVaZjF+cTFexU3
423jgA45G1BC/h7LGknXgKBh95C9771mO2mSrw3cW/1qP0ern7NoXkuXTPmc4LRMUo2MJ4y6hyBe
alh192M4VJnMXMQbhwiR/2jS2vXN70NdR411pMASUah4uhxWPTdimFNX0sHe2rshJZUyLXaxNL2W
RKxaa4YjAH+Pedfx+OS9zVV6ZxBNd3698ct6S5juwLmfelzhzwaFKN2SSMaDCL4+u9MUWrnvW7bs
qdo2VPKJuZTQXrju+B3LPAyHMvEqXstYs7KdaXWdsbTg6JYOTEai6s/fIUV0KSI+WQyQ2Oo3Qrh9
j2I+YurXjG3aqX9dWT0Ifk2rBoiNBnwGhcGI30zvDlzNUyElM/IkMGzXt+eFPCIOJ1LmAeuZVWvA
hCN/3XREeVxWr43kPVBOr5Emy/KNs1+BmaRN0aGP1MOM2y4ATPlZ/At2X6SXjJpjOG1SRtcdzlKd
NYdrF+KKWylBLTt8dZuuzE/tPvktPy4nNYKPI71pLize9Tpvilwh1/tViO+Rd6cOqcpPNaXwFlDo
MhwrhYk3ZvAE5xJC82k/hjJNz37QlX6Wvip+TmkJUg7UYZ78OATwUl6xEPexnQTLe709XRHlpo5/
/ytEwcwZXznlpEkdtVl4mGxZf22HiT+y3u8v3TyVtmtqH3tohdb9tB1Fba30WdU/gXWKy6K491Wu
ObI9EfE9Riw7MhV9MVsP65shN67DfXJAR5ofmhK9gj4lxtlSyJX6uvj+hjVGhvG8/LwnH1tyNVLq
L7Cy2XnORQwaZ2ETcaF5Vlz0dcGABMVMbbgF37kIRWPbCUrZEveUzlJm5shV3l3JC5nkNWDFtgTI
i4gM1qjn+OTaN2xH1H1ksu+y5Z1mkN5CRFbf7lVhO0DGcwR2vP4yoRlFzqW7ROTQHmpexy8oxFn0
eRze2nMqcKaj2qY7TU8UitdXDyEZmDrT7adUlSFwdqWCjoHf7GcCmToRN0aNfyeNi0K8OKrQvwnF
X18Na7YTESI9InwZqFNMo9M1I7LhPpHgXrpo2k1Qcg7xZptPl2kOy0/44XYvfkQd2fUJ/VqJO3hH
+CqeExaPbboWQz145h7lhhareFQRVzhriaxG5VcS0hWGawwpNBQXanAij34IBkh0zJOIkvslbcok
sINbfynGLwlrBngrvec/6OAKg60JIpFGE+s9IP8j/4d3qsruhoXqlo/OBYaKytRwqNT0BPPmaWLM
UIIkpJnqx9yFqWXwEsfhm+6PMyYVtIplhoO9t/wodQJkW8nh2Ij00rNupB0bP8T24fhddVis5gBL
hs5OPG2dWou3MM39qHBSmX+zddvI/uDB8Uu3BqhvVbAR/x/0tPVl67ymKKGo5dkkSEv1hNRaJwqn
L8vAkwFu1NJGtvhPKB8BU8aqlhlqjOU03pk9rWcgcrHkDa5ZFiIFji8y8Op0uUlCwU38Blk9ceyH
LZ+QrUHtWjxg9OQMC1NGfPKhUhcMTaWlxUhl9xbhv97CMYJ5NyG7GPJMIE2bL0G2QMj+1JbjNNIq
6eJLM86cv7rUr2z8YU45wJCipfJBl0rd6Tqm4i4VJfOB2yMiLjQ2oxsH4sGbneVj/zCAj2w2OIYa
t+hgqeTjUKTfcMmdIq5NDJs0qr39biK2JXsuj6XewvzoxGaWZ93Wts4FAak16CZrVNOvguqKSZ+H
GT4sS7pzF8cvzRfqr/IsGh7VODZpx7TT/W3++r8tW70e/6plBww0MdC3gXTh/Glwo7+BYV8gm99Y
CZccJaWeGUDy1uMtqYAaS5V7EYm0cWtca4aZyLgh+eBxhKoCA9Gf3GDR3xfMr4GZN+pi3oJD57Wh
s+xyKhTY2TBOHpeR1ucnfRyj3B0x4zBSdmyAO4kIbJUNyn/t9MoCcmU39nbWHjYF/52VCf9Z0yh/
2olsBlIUNrz2c1Xsf4NNvIpsYaC/3AGPPE8zEjeceBQrifsJpcvYd1KHinig60C/vs4f2Q02mFdG
DdfiBjC4EXZCYhxO6PpkMp9MFqoZh1fNLXlPx3rsM7vbenZ1rLTH1/Pa+TwQyo7sboRaF1/L/G6c
aF1IvzVrsFP97YY+1efvOoxJahsOVfSJpvxovZlChHyuzK8MMUlwu3Iau3O2zNQT2hNZw7txW3a/
PWf/y42smoAHZN72vCtrQewGW+8V4nKjIfyYYXwHz+xzw1G2I63dmXjbLycgJJ+y8USQqZPhkMc8
5sneMuWPaF/sUtREVrFTvalgmXmiOvp2m9uUelikHwMnjlcB6Cq1LR+7MKG0gP1b69p/frdt/K3+
fVIdOFRYuYAEP6zQAWkuayyPnQummH9ozqmzH6dR0He7S9Z63Ra3rZOZrU3T2l+Ms2LvtRCOgzzN
eug4yks1dnT1p+6+j1oA+3RBdQQjCJYMm/xrFgHG+Qgd+KxbFskud3Jpipc4adue29RVeRgN/VvR
knjAbYuAR/xeswC4bl2j92zFV9Yskm3tajwTB4WlG1sTIhF0v5KnaXcJzzGNqVGpwDobCosbTxsf
v1u3oJMHRACXNAD7l0+w2e7SlX5pHqJqNnth12crqgCaQ07tlsGNwjemP+cfdkttbElw/CGdvhym
+3uab+zDrqlvVf6ovQ6pNeiLXZyu8BeXsRhHxj25u9pRTke4qatG7f0nvMVCL2LMwBHgDHrEz7Az
mjN5/QljVTRmfNUaLKYornn6dy5t2iGKopUvZ688OweVQiKdaaZwhkjly4Y5lHXeoKz1zrDDWk/M
IKmkvCiPLLfyIolifHEi1MgxRcYezQ3367TQO5MUygReRJ1yW/z5aXY89dGENLOUORL0nQYHdjDA
tlKjsbRFOXG3B6foDqVb/L0C2XuMHvBttxLyoVPIMraqisybGWa8TjVE541ye7kHMT0aX0pW4zgP
p771Ote1npWfCA54WJA92xVu1FIfNJxTR/SB+cRQLTuar3d+NBGyg+NSUIcutSC3udTNWm0O/vEL
D3Pc1lqkXO3jeLt0wL26QhpRtlTYCiu875Vqk6HG4NJXtl9x5tNCR0MrESp8cIYhry3vb7x4UK58
h+xsMf4Eq7bK7jY2V3+h4ZXhqZp2NSpIQ/pcS29QVO2Y7TgzQuGtjEQ8pgyO47xL8B+lg3Cuxp8I
92sn/NgMFtcZTkWTBi/DOVkODJX9P0hSSluT6/cFH1rpQHd+D4DGIPvYr1QB7xwCLxjqXclRuD4r
C9jC959Apz1PiCwvGrZkqFNVYSBb4fTg5P7pyKssYHdgu5XF1kMIaJb45SNQWp5JkhXfLtd+yznA
6U5zv6dfLTEuGuoH4kJezBYgBTP7QJ4oB6g2VjIkZu8VrjKAgGUBWntWf86jLxCyFMVwuY59SNG2
iJC7j9rWbxwerMaMOgcR0Pu6P0+gRBdt2rXN0E5lSvfDtfJBwJX2mZzkJU7F7QAm0sWbVNwpY+6M
9KC2MYTlQZQ3HJWKCNCoZVSit9V1li/hKpn/z3wFkkldl3dzoBz6/uVyFEv1/vTiUMzDJy7vtLUg
YiAhnoXQY60r6A26nJ2KBoz+9ei1Ebi+0x61GocNNF/lxYyIhel9CdK+G3FyEN8wtfbjqV6Oe8uZ
6ThnFOo94KUfHgsw7gLqBpPf3lYLuX3jH0MmGtMwjj4WHt6FO0HlaTleN0/6RsR93/ZEB5KdCG4p
WL/9OwSasP1rgm8AkWXOwXlGg2j93wwyL20XsyXmigxLdpYkFnp9twVmlfVhWatBkAoVVdEHoT2K
c/P7puLmdhnUbzRQBeHIzZAPyhasHAgE13ZH7k8bo8oR6MgsyJ4H8qJ0m/DsXgIBM/BmCw9lKR0p
Zlc8vHGA4Wsp+U2srwnHEF6IBoaBFrffhSobSVKlz01tg/GZNkHcBooppOAUhfiUvV0ZtTubWROY
1f2er0Is94bzYshTAAUbWtS4XA8Ibsv98/qTwV+qLAAGsdiBnLu4jC1f0MHukLSPJkaZFdjAmwHw
S9zPWzCVsDNurIfOQlLilH9pBqvlPssJQ2SCWARwl1YMQqAzDl1ypPNzCAdo1Oz1pbF3a0brvc0H
zHyiYH18Mzghl2Xc0HjpdIAthAbE9s9uYHwcowuLJUVclMT8XaVTQB6tUI6fwXl6qiQTWr3R0sql
ojSgFuwMkkjfLMGEPu8c+DpId/OFIr23XaHgpJrXQe8bhtPYj3/UAjr7ZFLKEoAZUYwTd5egTmYb
bTSks6YebSxvlpfMOcn6G1Z+2FyBNP+nGhfGyc3kyLsqqKmSNl7mNRZBIckBxAfOHfqBntvggdE+
ULExqxRvv79v/y5DJU2RV2vWhaB/9kJN0JR1psc+6szP5bFxHHAVHbt2XwGERCNVxxMq+/kAj4e9
GcuXTstLfzKWeTYJhYc+bXmvtBYOPO+zhLbCeCse1LZ5f49L0yuZVQbVWBHKg4cE6+CklqgdJcwa
eiYVP2mIkKB/sNILyabAx6V00jw0il3VjD7J99NXTTN/JQ3LgZljJyemC/c6MekMIgR8/8aE+k+R
rbDBJf4ry+b8Y//ytMug+nZMI9Sn6+hGT58EMoCZGKi9RZE74/EGzAzSIqKSNeKAmy3OMfFAwXcy
FNYxzHQjPiUYRYZzUlYcK55AKAvPN/FL7h1qW65EHNpxESShO3uoXjjpYdpXzf1ERJM+KMJ8lsew
Pijk07rPK6pcksmYvDbUfRfeOBM8rsX+JXLmhZ+vVcUEN3EM4M+SWNk1a3xgTJRUe9XWTQ+RwskE
cmsIjqXGA01RvNWUo3dWrp87PGGYLuIf9RMMXoZF6n2jkOAdC9KOWbBea9+qqnpoREz90xPg9d+V
uxpl4PbsiRV8qjG1KPRAHSMv09mZB5NvRTjVgAszyDEZ4EmbGC6qpD0fZstLTgBLlkDcnu7Lm0sm
BY1Cq75oah9zHrMwzpr8avkVtavU+mSw54+K9fgsc02lbkJPLyYHSnlFitofO4FCJE/NwyPQ/L1r
zxYcciKIiDzUUz2gIPstogXE8NgMqE5VJnHl1ivO88GNHxk6aWrbJDkigZqHwulWpwl9282d4Bmw
FoVR1TsdKLQ/K2UB/2Fe42b1ihzeVdA3HjIWUMFddKYyIfqHrDqEhF95fYKAMPQU7z0IRKokMhdv
70GiN0MQPrsnZZFbKcbYxDWlXJRKKp1Cy/H6335uX1YnIQLTta/HRMsPsecNPZ7fFIK3ZNwfCLYp
vXITWxrDt+xnTkooEJuffDWfvmWPP91EwrUj75CFwnuGv9gks9OVzI5OfLW1fWsovcr3S9FTTqoi
7YiW1bmmXLAB0nmq5KWZqNMN1dSL9H42u73syqdQ/0dDwbfycRfWOixB0ejj1JCfbVNMWAR6qpQo
x+X3cyO2iX2TJ8TdtxeohclJ/yYnappjEGu1TTVOp4GbNE2+g6ZmiUxnEJAIoNRmMvpZT3Gy2jb0
t59HDp5xyJSJ2NaxcIY11J3gwM+BI00Om97RuXGOxq3RZsOcnNNyHISOELWHIVk4wpU8qvB6P+3t
vrFJGeLQ/3pOWe6oJrZyo5Ty5fqPrxDHSNdcgCfuLC1RVyMrEv7KvqcOF3XoMTFCG8SKupFRHPQj
utMCS1Jg6OPHOaZvtyu+kvETVlczwj1hCtBM+pOwCIZjJcCL8QCXnKqw6BvWkdVMyKK1VSesRYrK
JKSisQa8Kb1Yvspq6Pa2NBNVW+X6HMMU5LHdx4uibF3kONT2ndYchtleLZgvZzwMCNmWcbwXrfU7
ImWYsc3vJFLeTk6pHsihxnBC0L76e0FP+kNpGfcqELtJ3oG0KYTJXLsil3GHdCSpfouZxTbBXw3n
X2lp/gAbXvPCzrd3yrLOKjQGjHeKQbENdP5tiq7dmEUoCa4VS+m4zBGiBKlhUdyWc44y9KUYNfnD
vSzoxkLVR1X3t1bx/M5WoxAR3iAkICuH84twFqWNyI5IG8tFssOM7peEbjgMiEIUVNiXJzcsJf9H
7M9L2Q0UydncoJzXkmqhRMWmzKCVvDG9ikt1ZJ2AG2yL6cwAv8qImb0nxxCtXEZZo800ES7BgV1W
cjDRRknjSPqTPJpYsjh37m/4vrOsjgci6NJxIzq07OwKWZtH7RrCnvO8AqKma0+yytUJWHentFGZ
Kd4zJNqgfXHgZIP/djPN5I5yrDYcYeV5J3PPgddYcfZ6JLqPSCeF54LUemKJ1oo10zhkqzoe7Q7V
1soMcPxcRa1v6ocnabWtVVICqXgACL6CbkRT/s6QkJCFnFQMkPi+YfVOvflcAvCz9qK/ihHZRFAW
1JKV/OoodT9FpGgLwyycHRb5iuTSke3PCk0xwWjAFY7f9kBP9qk58uly4xRBgwr0gYx4z5Xsab1N
vL13+6NuQoH8bIbPhjj74rUtaMw3OQEtt5EHq/JSslokQDWGADHot9IW7iKtbhKuC0summjYl2t9
0CDMwVTbeGUszylOVy0eZQTc8m3pSbk5+L8XRS6S+qmKhk54lUMkXMNoVAtI0PsOuXM+O1uvPwRm
0t5dTive6dQzzoY65CtIt2DlFlNEb9B2ZIlkhUr+SxK9wBUqMrpS2GObFRs8sx87aRyIELaz39YK
yewmmYoAr3TGmpZuW76dk3vvJTSmf579xcwOzuysxeO86dUS4iPVsipCPXjwGlT7m2OLmQqBTrg+
J7Q9nkwiykRpdRnCms3TX5mX0Ysyg5OyzTFpO338bRPWpdgJje+Y3qqKKgtxUNAeTpYyn6K8YUa4
GBHG0mfJFRPuYErvodxYvM0Y6HK+SPG1cjYIjsQJjEpaGVnP7sPpe2kkUQ1yaAaM8sPku5iCBemB
YQfC0Z5FY2vTrf2f//C79wbAU1+d5boneWD6zTGwmghL/A/CzSPGm7eUYNJOyLuuC2umsB9g4Bqz
GxRohCqkBZLjfaSbsjlg7BGkfonjrfDtbMIYPwVqFZqVhnY0bEPzmSRIHJLo8PmYqBhJf+yKsYIu
xFZh7+6V3sRnIOuRB6UBrCj9pLW41rkGWv9Gb01YUGgbE0jg6iYidp+6U9YC+xCaFOx3xClmCLxf
5DFFjJ4TPvcQNYG8Ti4xL7kRdz+D4Thd036KBrgoh2GVf+6bvAj3EIOC4STnqpZK6pW0nAf/8Gj6
GVYdA/Hw3d2T8ByoxknHe6mTAtLK76NS0oO9k2ecIXHnUXnrqDIXD6A249tQRAs6EM82j1sAxRQJ
j1PTagPsYtVLzLtnqF93KdLnYV/dRzcjEVR3gduVV8cZb3SWeLRvzUerFu69NQqQ5G7bYwMrLKdW
kuwPTzBHF1dnCoJxXCYNp47Awz1cif2640jIMiXF2OjOdpAI2hYCKYbxRYrKtHVCmXjwUEiGQ3/4
G0hF7fKRDqyGRSLNiX2h/0nnu5rWCJb+mOdjQChAJ0M8kUEvEhXXEar3SZ5iuo91b7ty01VBrDWj
SSYFcN7zG0lQwCi9cQxKxEb4Lk/s9zSkGV2iOKKIii5TAGRNlQooeABzV7Uo/IWhjVweqUjGpUsO
fWPpLowLCA2Upif19eCr0gvCW6auo+UE39VtJIEF/k4m3rSSSsTF+nbsZhxiUPWu6AQV7aOsplNo
UKW8XIsd8q58oShxnQ5UbkIL3qz6hppWciIrmcBzQJrj0ySxwUb178ntnUIL0BQNw6E8Ps9VMzOy
/EKVAY4GrkHnTAxYe4pPg/4iY/jw6WYZNZQcwnDR9t2G/v3Y45nNTTpsGR8byphJP5RnsVTHbVv0
ER6lj69w8PrYRKRybxhlW2UZWBiz1BccvgnWiqcLIM8PsusiCyQjCgIOEOIVaN8FAPcuvJMPGnNO
hg/aieBnJiuFQxLfaeXfCwHRNvizj1Mf+kDPTRnRNh5ppyK2XLOw0b7i9NtSsBUc+yVZmeFWIlhF
1+2Densi4dmx81Wa6LspHNGDKvxA1PPrOS/JRYshgQf8o/drmbF6M+gKo8Db11SCBGu965iJhW3G
0qpHygqKJjmXCgKgiy1C2wA2drXfVkPbOQMhuZPgSf3p7cnLnBWcXkFFgV/8zwzpMMuX2paN2Lou
Lg7+TwqwgsidSOO8ShdUBNw269kwQ2qcSGw4xmqanVqgE0oEmaJWvNmYLOsFqOyhwXXeZNULgJ7G
e04o68pshzIvFrn9GiB7+gf6WvajXDXCQHqm/5dltZKX+98vqodhl63/XAde42RpH2kxBlOH22w9
/V4m3ihsZzxrD/X8GCdP3ODgwPkr0sbblhVhqFr29s58vFyu+tnjXehqUYgoxau9tsMfWgpcc3sp
mBqIU360rOm78LzgcYGAqi/7kOwllKhhaeBDLH3Q4LAlXX9IodpaAaWu4gCL8XNLYDF1u7Zs4Q99
316bFakv9rwuMHfapE2xNR8YWz+NkP4+2ve+aoFyfdQavYGDVR03XsTGuoP//HwFLAz9xRmvLQEp
4W3gncK53cYYfdtQfbM/EjPqxMXnyHLrt2KCLgcLbr792NOs+r2IX8lZdKMLQ0tPnavPhYuIVrtY
CpUG+J8mmPgSarBkXFnHgKu7YH6MHxqm7S2dwDRmZy/KJOZ0x1WX5kcO0qknN1eaEA5EQdKazb+u
lZPD3iYRJRT8o9AKvnYH5nPW11ABT1d4IX9RIXTTYQg75K0BhLaR1XkCx2H6aFhLGwJX8+haouaO
h2j3kDyMWATbe3tW4hydAqmdYjCXLcx4rvD1Rxneg34nw+qbzs4aFnnsc7YrOhZt9fUDn4RrBK0K
uZ2wP+BrCL6O780brEEWDlcOVpvfN5LeHP/KTrIvt6zoi5fonHc5WL6SPbWVp4YOzdZqb5cdduq4
nOrTk4tLxntLgg+vUBiZNSPIt8rW5oCnfKBE/SIwg1wUmsFIDuNGTX3Y+hnOd1ONBS68TQX07DNX
jUsVUl1B1+IQP9tBQpNXscxIYFvBsQJmNak5yiFhgbbnFqtpwnzPMUX6snWzdDrOZuxGCqCtIvK/
h+yLcFJlfwgd4aFLYK87wEVvnH7aFQjlVXhkfZ9ylvHMo2NcyFZPJyC4exZ8yWboOZ9J1V2/VfBA
1VLH1aEgZyVTAnmbznofCKoHIG3dQu4RKvoHH2BvS3Oq3nt8Fa5BQmkR0/0194hn+Tl77/53j1el
vOva+v3Ik8RBcVgcaIjtM+D8MeaIQy1yE8h/ESz7nNZfuQ/nDaxwqKpZ71wVWAdsBS8wS0fqnkmy
nfnsCqrXyzXI3TZRAmuRNyHHZbVW7Rkf2WpR0R5TnAIIpiRjIUkD5S0J/OJ4OHlaU33Kb468CwXW
Q6YUCro2Sq0eDYUNIaekpP9a7nl7HFaNjRIqD8YT2DJlCInwbcY9hI53pZeEMo+cjPC3ph3TLNGF
jiZmOGdygOP1ltV96P8kkG5pZptuUz5bqksgda7MQheXYX/AokfXnQ6q0ZAn3+95wWXv7yQvoCOi
K7fyyw1ytv4KRhWlkXzP/AUTRhGJx4GFXDkMyLpUArmSKcTRSm7E8qJta9LnRsdg9Cc609uAt7VE
g16hg11ECTyXwEqRqSiwqf8QmCkDqE0xTIv44gFbi1erUrghVVWMhr2E1sclcv66rwOlw+vlRhHd
mkiwox2KV4s5bmRIqAfCIrAmGMk8tGqlQuTueGXT+tpKxM16r9dlctzLexVWoQ6wmCzBcA/lU9Li
N8uIaY5rhTX0AgLbj0zULPgeZ1yqc8LBBJFN0eydYaW4CSz2BSCDPrEvuuzPZAE5OaucKSiS0Upc
glc7EB7BFi85uyi653axIEvOcVgw/lXTx0HEFPZltQla9fJQbOZI/Yi6t20WbOD4DwfIDqE3khKD
Q29RQP4ldOTGKkp+ejaVv/0S63d7pp3x7kleSy0gRFmcfVImuyvdB0c/SZ2G95jV+PYYQxmqXd8h
fZHXojsZDf0GXMdTbWV3JUFitOjJcuWZnfL0xGCAhTFVIcfAuqjCoU0DR0UW7Wwx0h5Pco+bZ7SF
E2JJ1JQ2f3kulIGHovPoS2bC8Dh5YA64FW5DlmBcNEj46YvitzDNq2qmb0T4vLlBIF6hikx88q69
vGT0hqcTbaPIYo+ZCJuiuoeS91qR7lDWCNqqG07cMBFFs8SjDZPnV0fwRz2NNMaViYYzB/Hp/tA0
9KZcwGXfqiyxVQ5tfs3d6esN7HdEYutHvzH08nqelSCy21zBDD96yMAyWRREpeuAo11Sodn9ZsJm
Ro7kUvXbhfMinhHZX6cgzP4ZQOK0XsKaqX5kwJuJoqBmP5YyeNxCYEi18OPKrIsA/0ZHaEb6wKTk
m4ZvM0qF07JDM4OjUJvSiRLve674gCI0/9dBj/2WoCA+Q+KCB2S13cACMCdlsJ7yUv+guq+m/ClX
uS/yCVAoCtOMUWSCXVuTfH90jFJyTdkOu9f32R1Gp4bbZ51TGtuHZiblzPucvc4qR04fW+aHyGvy
/KJws5UAvpqORrf0tI2sMPE7Ty3jLaDC3MDV0JvYlJ+BEr0LWoTS9hx4CikOQsny6/aUSDOQptk4
U1tdy5nfBHtZOuktUe+GeCisbpW9/FlGy5REyhKmlEYF2nQtSWVqpdz7ZaETBAS89DOeOC/rHGfp
NnJElr3BUWUzXerD2PNv6W+ETE6IYezp2kFsTr4FkEWdLBlBpoIvEeZEhLmIH6GXgW/1cB12L7n5
rcXUHnxsmmKu/fNrQzk/NtoKYo7BXysU+Y3eVqZWrnBGR4gIModRRSqhYVJe+OGGvLgJhBauD7/U
g4rhdeGim2cuAVj32XM1xFzY3HL0356bCiObG/nl6qYbVYGfR21OM69N2IH8HhIU7NmjBKcNM7KL
COeN9V7rLmlgKEmWp7411EgeZBbO6shQJAfld+wl3qX0DHbB/W3mez7Kv/9SrNj3MdEykYGrzcNp
qFJ+ySrFRoQ86DWbicd36BIxM5zCstoIMrhfg/WnR44wcpwiuRVYbKChv/CnSi3P9KIlkvYl/l+3
ebYWwLIOoAUcxdIlQSOS9B+wfgdGODGDC0+6ORc8acnlL4tRhzqvbvMoMFRcIOJf+8C4KEJoobGi
85KkfAnJnou0xPcJK89pWbgMSlo6RuqcOFPpXCntNLZAz+XIdcWqayGDicCTMjFHQsyJhkzVRI/D
7n5YdJsElfXcu43FYf2+EEgMdEat6FBx15NoIsnbXuM7Ib1sgj47kLDEX+r5u123g2kkoUWoQZHF
bUSgKdi9B3qKcEk8c2dwjpCJMx13FKBJ4TQo1x/hw+yU+k8+Ls6GBQ2IrV8KfeA0K3UHzfXrLR3X
HaAJ3NMSRqC/AlJEASqiYuRHxIt473RfJLffGS1FXsfUZp8abH5C6mzsgOjWZVSw0TLfUjcLTJBK
Nl2K7QM0SR++7e145E7GGYG42CZO5PGzu3/t+0ezrwxztYF87ZUCGJ0swYwu0UsbqJwG1wnsD9MQ
EnK1HEKbCb7mfUlpBXav6pBgBBX+PYtDyBiYC5mR5VHfWECqyYjEbbPzke5FfG7UJy8qViVfVhsF
EBaAtHQtpqWBu8QxwMfIrAOysSdaI+x8m9/+LidWxf46NHpE/YPJ6v9ZEwTnYZ19luTcKnQE8JCf
qP02jJ2G5bKTab8XOgQ8gscxl5j4fJ+vzAnwQ63P4pDLvyu82zthDGv8YYseU4ge69bJxoNtG4DJ
baUq++eEWGjfRUORTPY6bpwcRk7riiL2oSTjxFqLzA+P4rXQ2AH5Dlg3nkDZg99c8kz+CSsHaIkm
1JP7+4jRzC9G6QrTm1Kl+0oQ/Ej5gqBRY5ZhliZ5ze7Cg4F6ghvA6XguJAF1Qr9qB1wsRLLj6YpM
YkV5RF4wgetWEMBoEkSujCEmXNmzTxVZwz64rK6aZH4YC7+4/AAKBSXHIrjsk0YRreRt+ncnImIF
gMoliEvMAcqpItTPfTRUn+w9nUjZnTnlfU8RhSdNU4vUw6jgWHs0qjQ3VhSiDIDfleNLgGkOujYj
pZwdOEEsh/GhYTa3j8pE9On0Hoi9sMotwR0mjQ6sxOQyMBWsIxmCClPu24Cj7t4qhsN7PZhYOpX9
mYosVHHwHZEJe2a9eEVBvWC06Z7qqpA/gwqAV1UIFN09+51fRV/tM3g125jZDcH/bUko6fx+Fjhm
O6ElyDBkhYvjG6jJ310Mj/T6mkVUI19jYjQI9Zr+03aCg8cHZNmnZWfOvGQ9UY6rner9pQYYwvlT
qHBTqsJmm2JqwXp0h9y43L8QmmC1Q9GmbPyZdyQG9vemG4O/ruCCMBn5wudg1+dBHMdOOc1MuJQc
WYAgkY+PfgfBMSLg6Lq4b9iimK4nqWV1o61bK/2IMmjKWUOHVOAvU/H70O7ZTtTc2sprJAN9FhGX
nCizSFzUYWgrY7oCI19HVlaaMc7Bkw9kr3XPmuz9CJC7bXzMUN/59LzcvPDYuruIU+ls6WhyDlLt
yOMuzhbJjILB6UF6qbRcp6zPl0leKsEpETYHBco1iOna5FojrErGBQDB3vcMY96g4vE5AGCHaLJz
PImFZF8GIiKvtYWFh6oIRQusu8ZD4uLlCC1gY7DroS2fHRJwcII3DqSW6nCPvyljyiOUjQ7QeZRj
KA0zRTZWTvtrzEMWrHryijyJy/RvC0Ktpu72rVhLAOVnbh1oMTKRT7Cul473eAjXltOIiCzxqUmD
iid21+6tMqKs4Jty6y5sEd4cimIf6xonIKp9rH9Oowd6ib37J5x2ulNrKhexa0LS0KGqkHJyIV/p
27OmX8n61+BSR/Cku5OdFvlGcZeNgKGYwWxT+Yq9yip/paCa9NiRoPtMqx1Xczzj35lGQHsHgjLU
1xVq+ts9/dCUb71/40Abi12EJA1SFu4P7t0KmDyX0htf7dpPs3zJgOeNt2Kzh7hEiFQq4HJg1cQP
c8Y6jCGnuHk6WTsyTPEVfZHP57vH8wGDkQa6XOsxgu1ej2lYUwkSVkQRFQVTtgEwzVpyYlVRBXzX
59awS6s6TnE+0gcLsyoDnX9KcyiuBn10HUs4myg1Cdsd9xFknujBF0N+2oS5ucJtXyEFpYRhX4Yl
rc9sa9fI5YZ2UBSKr+Yl4Lt7787Pevqq8TJI15Qe2UD+Uxzf/IFBmpYcbXJy1Amt0+9QFiXOyfEU
7NGCasEkX96jic2r8sORcos+lsf2LitU0Lckg3rVu/4pIUvgG12DwWY9beV4PJ/eew7hcH3AKiY0
bgimijNe/yBdIXlCVryKeWg/o1p2523TBxBvfo/3KARvL7QcYopwbRIG/xS1sNTKxYZtLJCeUy0S
hOu7JTiUHYUhe/IkfYYAS8raTrUkn93Sx1omEewmfQmCspUerwEdh5zPJz96ex8Rh2yoZE+OOPVZ
9SgALhwqUiDMkyxOO6cpV+9BwrWrpQ+xUHldBYtr9TOzP+ANhi4qfLB6SKmOWL3ShC6I8FcnD0It
c0EawzPUmr3tOSgFAGG/MGsd8esMRhP0Drxz+BCqfDyKVfA/C5+2TAuToScg6ohxUNt6iJwuFHOG
OLRiARBB5ImNlNpSnyMrN7e0nXGGoOVjPAqr3BqyfqZDi7RsKXJ9Aet9u1wKdbhn1erEX1amN1QT
XtDu7h1YgCOBSnRswd/qiALf8hJ4nuTWmCt1P0jfKJU7zSOGSpndfGalxAMHuhz02/+J5GayvOMq
Qo8hLQ+y7mdWKuhDDieT/S5dMaArU7bCYI3zOWgBc9ldUcs90jV7k3IPuV0iuEBQTtfRtn3aM5Zs
FYqhSN+xQO+UVYM20dWGxeOG0D73+vV0Py82WtXMEvJgfdlhPZPjoqD+4bdWkSX9BW16g8Ikdqay
8Nvl97O9711EDlDhYw3cyetKjHFlEr0Tiw6yb2nmjRxOCDzd8ErH+Fy92U4kX4GU6Dy0mqaEfhGn
dvjKK2sZIKfsv9v+9E2bFsUzDB/rxtCxHCFonmUjBQlEzMn6LMfd7h1YFuFTDurZPBWN1RdKOR19
OOAmgrdpFh1SRzkEDzuBKR/8xyrI6WX/VXG6CuDSuA/uAKq8ogBk9qpBKTAjg4sPye6/hTXF4a+v
1TUCm640kKPz2OPKGwmUvIsFQlh0hM81dGmW93ry43aJvpCF0pCSgkOqEmxwsZB04ZlJPiJOeWSR
gP5fu7iZ4o2dj1mM7/crq+9DWuxXF8wbjIQcKSWdDEQmEr0dLSx2q60eiS5dsKmR92XqK6MsV9Y7
tS8EVElmLKm2w/J/5mLLS8qHC2/AfvF7D/OPO73MO5mZ9dvrc7nAYUi2A5gsVj+xfrh3oMEWNoWW
NKZoGioVyjsKdgbY8SebqPApP9iX0idrFeUfklrO6wwj48AP86HOU8ONdnetxiQRfIhqLTfJEFyD
E0dBKXL4Q3BQFaJxx0F4zE1InnblRNido1+vipFCDKpj8PrDtnINMtUvyKITEKukMNj8pu598uu2
AY+8T4IOSl1i3RhGlNjs8RF5OICryNukiDcgIi560U8r6SuatTnhax6sANTPFZtlhweKYdB1RjhA
L2OUfavRNadkLHrRZMVGEESSUepdbe5xEcrPk3DP46khpIV4wLbGq0WrJLYCxcymGimDb3HG2hXW
YwIkBO/zciSfmbTgDX05NSMcvYOQ94MkmHkTBCkyYJ0GOQkFJaRoMi/Qi7RVql6K3dGbzIyJ9BwR
QOxODiRi4ceHKe2wqzXKvFBkgDePGV9YYixD6aopLnnKxR/I3m/+2ZdtzNTTsqpTm0OpC/kHalvK
SC9Wm961KGIwA91CtuZqArV8Dr/Aaj8D7Ka9QAj19vT5u453ospvR7zTMEhNsJDWlomQgqFubogY
3AHiQ4O1IJLwEiU8167paGcxEfJL2g9uN9KWPy/PXQrh4v9b8cq+9urT29zEinxw6nB/+UgEMY4o
lYvYOumLwehT3LqExYgX+xpBEdBUZwtwW+2TEce6yLqCBeQYCcsvG9kRGtRqd3CIMgyvCIuhNXcB
iDGPnKLBZaK+GGqtxjq4BX8hS+fBAyIeV1HNJErJGoMkwMKgiBjeQuO7jk6ZmICsrcmbknZFGwcO
e8ONL437A7zZe8nGPSnaN65I2X0tRYgsbdJB4X+Ncgugn1hjdyqvdQOYXjkZ40WPWxx8vEK7FObg
1lgGVoxC3CKq5hQzwU8W3cZ9xB4xrGRCKnTezARz+u03h3/Hl5NkqQdFognhvUnreA+0r68kU5w1
eXkBTx6oou/eEWxaF/PinRGIYU8drs7q58JrT55BoNNeTbLqMMVv24ewPdbioRRHv5hYNtjixwCi
833RWH7MSayR3ar1ToXVP+ykbUpXvRgVNYll2JK9FHTgWlBF8ofWOs1pDculoWDnH4ISz9PyL2a6
nZmUR8kdI//OQe/D5UxyJZSC7jpSnlvi0YvAFL1+cgrjd3+/4icqinO1wFddciqlL6kUrJEeXSQL
UVE8x5WQLry90DCGVAlVwKKtESo/V4MPw1hX2qMhuK9m1sldAKB3Txgjs65sNKwjYItzzQPTIhUs
/gD/Z/JvrK7zqZQ5ViLBoRSHaY4HQlG/9YgWYd+roGLwQU/dzFgouMKOG1AF8CirRNj0iiwMr8qb
hJt0m323VgThwU1QDdxrSMwCdXARNFIFsU0Tuzag1pGW8E81y57vgVDJ2UvujXdjI5CoGPbRegB7
FzV8MtCf+ShAOc+0Jhzvvf1teJot5/hnZyTQcwtnRYhHoTFBMn16uGIemX8GPjNOyNYCdK/Qro4V
Cg0wLpB0/umlDRv5fTcZ2Evga6LZ9E2SgkK1uzXbn0yNVADgMaMb0q78Txgh4WdQOFZXhnlqFSXz
7ob/mJzRcTJp6ACsQ4zuZNQdCkJvQhM+yV8ydoihoZE6sLxTLa2j8DoONMbWiEZgrli41Z0r26pR
JgSzglWvusNT55gCquRDngdtJGdyNL6YCM6TBPnbI1DJw2wxBqUIaSDlOE9xohG8XhMzmrb67Y0q
pSGq55l183vkoefOsqi6+dpgeFHjsU5mwqRvyL8tyi8eTUW6WbZs7+t34w4NYf9wQAGN1jKeV12U
/jjvc1+QlWIEBe/rObwY7//xQfcNG9PFCvGlmn42GfapkOe7Ptu7gVMfkohkVyQBEXtbuz91PGGV
ZGYLEpVDhsrD4AKfPLWt2vppEat7M90BEyasqZ0EkWv6+ndw/JmSGVp4vUbkDRorBeAjqqjid4lV
WERTbFCH1jV6ca+kAWUgCbe05gefrlKUKA0lc4McJaZOKdHkg+xedive3WN4xPMj6fj6hRcZ4Z46
j+GrLa8/ntA1xJ89w00R2iSmLGTkZCoBHm4cDmNe+xUxM9luVaYjWiu07BNKzE3sxlXiYq4ZeTFF
T59grNQ/5vRvzfCvpqt1WnuEcpjvvw2/d8ZjqciiD9sJLWpYHtswiv0gQJLkZFO8YZ+L5SYSV0on
YeSfb15CalYT04mewloKyCf84Q8zmulFkswjp/3QlHPslaYfqOCsilBEskqrulr+O3isJXEx3Xt6
0BqIa+aJxp2mCPZXxI9rbLUgX6Khr9qQmeYllgrW14ri0OO6AY+WUJ0TB0tFP3BpxZv/O9PxPh1u
HMQ7drbY5uAvuv6CpOIyOWwMGeNn5MqkVHJ9PsLukPTcaKOo2LdpuYSJ2CMi9PA6MnILZwJPlDTl
o0wQbivGdpWG4GVz/5zDWmniFsV6BepE9h2gLjbiUayvSXHamCLANg3Id2AQFr76BBs5b2MYD3Jz
AGKjH1vWtax4jkhXoxnwF7jc7JUQ2wlRsKQE+FZJJGlb4BTQSnZkvIPbP1Genmyzu5VzXE+aOa9b
p6YEukbvwl4qe23tGrDbjLn7QItbymJfOcUYRzVds2cgtyyUZLiLmsngRCsKt0iPQMrYo42dgIBW
vU79m36SlGCQJDPHvyGj8L/IppGGPgZCYTzt0OfZWnWu0NmGCkuBITuAF8j0XjGxRThaS8gUlSuS
DX4qRVuXgCZmL3S2POSpxRpazZiOWjYfY1mz6bddDWRwy4CTEqzAoJg66MJhctFHrz72JLfIw8JX
NONRicg/OuZdEL2u3GprvBuB80/vKA//ERqcOwg6pM/C4GGZdAQ62bIQQW3IXfMi86AjS61uPgl4
WMBydlrjYHHy4ok+jKRnfYG/a7EJKDdhD56I7iPPMexp/s5W7o8GTLuo4DJqkdW7MbahWMFWkVad
xr4Zru/ggB+RDhauqdVR219WPu6j0Txp8FmJqSmamYxniXbMkuMkgIAgrAGvJjtgap/BPETbP00U
GKcGyRYDxFelFdH8zmb75p3t3JA3eFw8T2hyDH/RNb4VTAOlcNsm7Qu/U7ae0XCeFu9feOOtkEm0
0+Ox2aP5xKeouJBaVf1X3+eX9A/4oFebGH4E+pqCMjaqXTb7CDtdn7pgMrx3SzUyPiGoNrYQBdvx
CJC0KVubEcoopfOlOyIc8OHqv5KEHFbWe6TwrCk7FhXHlT26SeL1Qa0zIHgET8cylSUix5fqyP7A
qQT1+S9isvOHxsBQNBI0xDF/mIXzLBsTDUEEayph1jVK0KGHO5va/DcM3ajYpPGSQtf5ofYxs3HJ
LeEcsyytyw21S5r+Ys50/9q2ng09hY0ZLYHaXCiKZxoQb87f3k0tVZhmnpFu6YnOfo3aW1+1sUjM
bTZNhve5V7hgRkzJJu0wjQ9j88dHZJAW1G/sU/hANth/fE5yi7djameIZRYT3v85aW/vFui1KYRm
3WWUscsCohRHGbiTB4RDh1qlYssDTzGAumJHd0hu5CRyl2byr4mmJUOZmrGKYMmwDDEYuln+ZX3V
/VRJoQ/CfzHmtF+DDUyfPj/kzBbrKwzesWnc2UFMsJ6de3YvjXxOgG4/wbYURw+dRrSYyYL+7BPx
5G8wzdxIVR8dBW3aoGIpqFMFuYmWGiTmNpnzmUFSb3kYkTl7xbiq2aIJMCd6GgeTf1fHfU63vc7n
wqxvNuhdWHxRN09saont8Hs7BLa1F1gnsRyB9VbCW86S7aEKv0QsxoE3hKc+uUPaxZZWS6Hez33e
jTGgQk+wImD6NlAuz/6cABHfjrAKC5yg4jvdF1Gjk7GkN1didSHQX/skhW2fxsk0U1AN9C/EgnkK
X+OGSl9EU9zPwGnaRH4W/O4rjbFxp4EZ0ZOURyulohH4DIvovxqYJe0nBI4lsqDOkn9ao0EgglxD
ZZxKF2fQyozsTcKij+KZ/n3Jf4E0pJ6QSRitBH57ObBrDYeX6n0UwOXSU+2fnqTJVxa1Sm1tGMOU
NCIY80zI0DKtWUsVJFBVQFy5g87pnyXe2AzVBNj47nSLZXJELUfDFl0WrTJTDvvFNWMWS/P3YUiE
Mq0HA5PBKF9P2YVaCBxKkVptl2c89CNMJLl/j21J13k5DfvAFpVB3e/5eipADkiWgsNUFayJZX42
wETO0RWvgdf9d7wHtVjkkn9FZXqbicuRbr8GOzgyCfbHQVcSNvVAPZfGvsIzP4Jc4GcqamlLVQeA
qEdlMELDnn8L0iHFW2RtwSKLS0ckwSE1bmfb2N3bcxzs4ooHRaxdOCQ93JU+NSq8aUEPp/nUWd8e
THMcU6go/TJmi4cz80pgyK07FfkS7FtYciKieLrVTtOfZPN8feXsj/RGKkSo/Wi46elmhlxd5AoU
yMQ8NXSs6PzBuGzU27roljuLRt1aeHWSc1LvFqWNp2PtbilQnKJs94TwmfpDhZdzre0Fzgei8ygB
I+uY0O7UZ+pDg8Eu0rzy4bDQYytQiKhXsseoVe8CQ7XVI+o6njeRr0DRZoa5H/u3KNTXA9mxrIXe
HvUqJQjwCNfX6+imMZhJH87HxqCMtb1OZQnF/cPXl7zIXLsTstByPGRAOkHsrP+/JEQFlsMPjjrP
92+Gzx1DvSk5fGAuGex8qW8jloGWueDm5Lll86GoVO1DChbPYeJJpeh5N5OwGJ/mu1vn4ycuia8Q
r+BwkxWsN2rIZeff8JlcgnYQBk9YDmeqL/lYE98507qD3TfavvN044vfOiFIN5RWFPMq8J8PeEk7
v8x7YGtXKZZHYeEYCf2eFWsCzY2TRnxCL26WwKkHEtrSHNaPk4ABEmtn+AcB1ZRPHTokugHZ4jcc
4Y8vHVfDXufcWCDIaktpS5k9LxR1LomtYXouyrVNivjbtrsC/nI93PvZ0UmX9o+bSWlRTzyFuamf
h6Ujk/Ls3l1JF03ds+/mtDS0knUUZ8XTfydhuRuqJtmgddli2BDxGM/q6nLuTizdxvC3sKhFPecV
7jg0gtGY4j6lWGlPWpoi81hFyzP1ZGFtY+Pj3ME+RgZgKBkOcctTQslr7Hb9b4TH+DKRrn933SK+
DtTZrNLmyZ2lZirX4olgJfWqFSfO5nLNoRPQk//84rlskvY40Ucx3fYR4ChJkHBHxNimxtYu/PLk
fwyxW6K1hWC7pyHZUEaOvVFx30ekCyMe1TwVQwUP8/YepiprTCIPlcx/0kZF2rN1ZOnnb+SIn+rw
IyLMKyhKPnBhznVNWJ7Mu3BptEYeyBDwBOTJtJJYYmA6MyiN6vCVQWK+5bDp9UQCqB63Pr2MdjFG
hgC9O0v8yN7E72oLh/6VAqHbDlOYisDNai5xDEp2GlfdsDgPbS6fFoebPKdEqEjfgyheoyex0qAX
+qeQ/SM/GkMYEEavBs/ueRxnbeuVRbODBTsNl9ki0AkJg0eW3ABuorRMPI4NnMUOvk3SKRFQUzeP
osb6Z0pwliEzhr2ubl0DjLGOXQg5L+diU7GRFdCAd2LOHzTfMpvl+GnwOfPjELugm5UwgMfJIIAQ
s+HX5KatbRh274OcRi9OEHqwdAlNKVBLYqWofUqVQYpW85CoUb0pqheGPf/a5NNgLYqZLLB926E/
AIXm4wI6zQwQD2mVGOnFlAl3oG8GXeffS/eMUJY1LcPZICzt8ll7FSVVyq9Jfki1MOG3ddezYYZJ
GBLsR/JJ2dpk4Ej34elwzRwAWhtc7Yyinnh4lbgvPKvnIaHgzenzvezgva0Tl+PuYNhiSK7bddTd
AkZ3IrUBryQbMP7tBpSTZ9GoOVt/w6Gw+zc16vn4xYjHF9y5YPLZcT7hu0jk4Wr630Y9yZxzpuVH
e9XlIuIYTG6ovslfB3r7j5fAKua6txAf9qPnkvvCyCJpgyhfXbfXzcmyIYZkEy8FcQ7EaltV/k7L
r3P5QS3Ea4qclEsgQUfCyRfeBUtqXhP+YcunxxpbvhR7luf0ZbBIF7w+Peti8ifwHfJA+pASDf/3
7O5c/z6uIUQE3woUSDdMy7cLfKPqiurVB1NzjCDO8PW9FeDD11R127acsmiXYOvio0zU0cmIAliW
Hm5oAFKk2YCbCQixL7TkQNnAH8ey46z4z+Jbba1pLEdAjxMcFjSuQAW3QMaGHqIglJN2BgUecrv6
vJyX02fKtzv4Y29bh7hzBFx6k5YOITqNOE8lNxbM+1D2DmZExRJdPqAwILY3i9Um1mAgsGklTtNb
qH/h+r4wO37BdRH543X+TLWT6ThyOBk1J5b0P45diFZMfai6L3g+LoVnY0FArdk5yN7Y6kKK7qlF
rQOSWJ8nC/5yal+75DaMaH2GzwWXmVJqa9XDJ0YOn90Lcg4azx2bf1sfB3uv9KkHr14cSqlqH+A+
Le9SsL8Fgo4lFr09cT0WxA4Jq11JDMKmIr8Q8LSDqAg6CseaNkJZsNoecu6egCk1bLv8O0Dd/r8W
Dqu5nR+LhqbfyAYePIUEs7fKe5uJ9szmIhNqHgk4VKBKBFYA2Gtm4yHKhdy9eTAEB22yfYWptoui
1Ae1JrixUBhMBBkgCZT20zeKBx+uaP+T1uTqBg4393kt4Nin+uOB6Bt9PeZTr1dgaZi/0RT83qPv
aZVOswfYZJN0Jy7sz8Ve6Gfop7y00pXKucSCO9PeIpck1dI1IumUnlzDf99tejJ1QUiY+AwQGSLE
wf0pQMS7aTJG2uNd62ExddffDxRZHpvRx5LOw/jFwrYFUPGxXxRCYy7OPQ8PcZ5RDmF6hNk9is87
lqoiwNNZ3CiSmT8OneWR2z2fpRlGfG2UPHNqLVnwLPcb7pVe40YTYX8c71G7dKi/sWzLSPSb4Zql
4QpIhvuMus5OS1wTYhkex9PpDPO0n0nc6sEjU37axpQY+wdwWDNTiNlxsbom4u+JvuDgQLGiEfJW
HyWn+O3xEJnNoZ0eu4JnvlOOee0mOX8xNUWusyDlYu9LduWcQwOf149G5K17y/Ps1THKaxmSj+QH
mkpX7VVv+qS+mgGjp/VaJ+8FupU5fRYzZCvwqB72j1wDAiMmwbuoiJ+HiqDHM7D77LRwc4qkfJ6E
p5fEiHc75n5LEYWA/a+nXFOcoqRMtwLr+XoEuWhOiaoBWJQB66URuRMKmE6UWrV5yaUNQffuPzsA
r5WJOlqpUiWji7Idok4WEoUxBuTeapoXMrpCo+EZ0WLnL9qoakdd/F2XeNwNMItqP1npMkl34pj1
xfsngYcuoziv8Tm3vBwy8rn0X1vf0A8TqutzY8fwJsOkKl+IR1RiMM2796gSY56kwZ4rAh+q3PyV
agonLkv8dXZLeKovrV8yUKz5wZU2TmaIEn1I6ezu5TlTWR08MIaPYONAAlsnLQ8Vp05y34rQRDnJ
9vyGWOLhhAglCpzVfAGnA4N08hu9e+iDqUYcWYRwjCkOjubQNYpx4NySwYPIFfuV7u/crCQ5z9Gs
xHwYzNwzALofat/xN2wb/PQFPkml621Q3DS45e+cPusFGptm90ajCtRqqmdB7ZctD6jH7tMrIpZ/
k/4bwrplA0Pd5HpKXxbtah0QBLF9F3uw/oUha9QvPknaPb5i0HlrDyx/VS71iJOE0kIOAyUTWlAi
TeEANSHslgS7I2P4ZzNxjjcjIfN+s/Tl96BOjFjLPNdQOmn0iPWf+sjWlIcBLgXba5TF0I1Q+3Dq
TOM+MhwRvrafaGDgvw96CfPsUgqgHWgVyLy3y09apCsB/lp3/+kQIUffeyU1le6Lpfsnfl5gVKXG
N2TJ/Fp7hh2/UFgz9PvSfnqk1VhAADo620G27zGKnmmzSk57gkmjg/z27CIjytA6RAsYN9UlFQJa
ZNmy9Oxj78oiSaApWTfBr9pxHvF5CuIjn1WYkB3AEpYxEo6qvVHCK1gzFWL3kBl0fhn4JjvV5j+w
Fn0lGS2rBR/atro+NW0eZjGhsOVR26x5ZLNnFOBuW6fyc55yd0v2rxV5ThWC6IkDO/Sr46GE/8H9
Ow4PW+WQy7sC9qS6t2ipISQaqS0HACPvGJmHAiVVT0UelXRgnXgXtTfBazQzlq+DgePALuANY4c+
7bbn5fY2+l8yUT3g3wLVAg0l8xso+fF6FpimPSTxxSsVx46kSmyt+RfXVr85NqLyiAgPtdhGqSRP
1bOtzt8H4pP07v+zW4De87NHKs8B1OkDn3xAV02mk3rsJilhmcg5mtZKS1sLe1rRs6HVe3DyX881
OzxwOcap2t9q74UYGaBtEsfIJbtqD9aB7BTl+LxQNXXqY85smbqNAbYWxPWaU884oWe/Bm/2KQ7Q
oYdYdiyRukatL3UL5CFjVGsdAVTk+zbsb4LylggJNEIA/9n51wX8eyO4LSDDS32Vw+helqVR3/N8
e4GIzaCt4rwy9yKV9nZb1noO2K7Pd3qmPK2aslSovXEeRDoh5+nI6Ic0PjERmsvkVvSd7Bityyy7
lGjRoyibbnm5w38xhmE5cRC4O46CTZPYy4ridMFR81pyqFfsJjD4QnuGwof+RlLICimfrYLCByDr
JY/H56esdkqn1jN3M6jJwM+t9G7ClAGS4U7fmdL1EU1/dm3FVPYMNy/5kWHHNy9xVVLeZ/JIh2Rk
nuky+PgR1CPpIjL49mSqAJ0kZy7yh0CUAnwXdNQ6I3CkBLl10ISw8MEqEKyelokaiiI0Bej/d16R
kYvQbhYkIMlY/v+oXKXBbpFl/2Xby1GAVQTf5W5bgXVDHdWBl4hEJzInv2W3cyom3GTyBBQrc0QV
oMJdHZzFME4pWffijz7Zn2C4/YSBIZsfo5uENQX/8BVv0MfpbNur1OhTr0vFDwe136KkzjDTnDf1
DcNvJ1RgI3g825nDIrZ0WWHExMOfHs9AVd4RROxLmqEyAy2IVNBYZeMe7aEaw2zvP+GyOjl+6nLn
1LVm7VazECK7RUAtl/OgByFtM6vu9l4e6Qa52Fy19XeBGnuVOI+kQmRRfLaIQrPvwVJSEkFg3MG+
ugu0eabV+lTCkwZ4kx25hXKKqIY6WAPnkXcrcVfUXedLWFey9anXS84AJStctbs7h7IjIx1aXFkN
cAWyFniyT0Ls4ui1lrB+oHt16LFLgXx2ExlosA3/vg65Aur65Y+ChQVvh3cRTKwLFgS50JIukwBd
vFxjMfTByXRODxL/tiKSU/jDMOw5a5r0A0fnUdNkuHpvEuDk9G/0Bmdeu8JstbWvCBKHDylH2ug4
/sED043LKbyNPmnmPZXYDahaWX03oUv8kUkVwgDipTncaAMnhQv3jfzG2G0gVRkG661G7Kc0CZsx
Vsvlq5rFlbWbQXzC6HdwPQ1acRbMzTYh9cQh3mmWW7P2G6o960UR91US2l3QTuKR6eMIKK8nF0aC
YS+JvY/PAP4wfKR1hPITZRcF//Cdj2hxWK7sz4e6IFC9U91+p4EMc5+6MZHNmHAK7yqX+j+DzTR9
DDGK0YMFP4a7Z6uCqiccxMd9WmFK+UAFqxbnZwgQP0I8YMoqu+OOeolH4o+24CI1h4DGyOKzSO4h
knCk+zwVL3JTc+/ReG2fJdT9wYDvHxYFVafrk28GnSPvx3u6lFl5oT6GA3dyV2budw+AcHVyPCR+
ZLX6ylghrS9U2F2Fz9VwXdTAUEmCkqkKoRZmtBMSoodIzSQvKn29WthvuinzSpC8489kkYdifhzA
gn0y7S9slRAMgvV97owOLGTsxDhe/9MhlyJnkA/Ut2rVdDNYrbYM1A1C9C1OzDZLJhC6BuOhkddr
yB4+tUhzmbuk8/PzqxyNdKznhHjS2/sTt/5fBn46fJFaxKg/1sgYKqoU/utX5dFatNRv72UfbnRv
3ojUZUpok2Fxx5xmqI9nKizODkBfcPoGodoAvLBtqQ2V2XiA6/XAAn841V3Iu30/nJm4fp/VZfOj
8r56hS3feA9V27bDoa44bGDi4SSFQcZO4i9+HWkiniSPIjn8yUSBBW6RMIulhAPqPrU0/YdS10Oh
/qNMBT2uyyUrqVWUzOQrIte6KaKXMzlQ3U+oTNm5j0TjGc+5zprlur+eql89+PST0f4A4XG059MB
Bo6G2wp/7neq/4pDI1a/J42aKQ+sA5XorMb+5js3NqWruMSSVcK9DiME1nwxiYzyLd0oO2xJ3uFJ
XpES5DgLomURUCOhNcqaSLay1Cb/kCEQ4mqoeHkBhqeWpFO84RzYXCl8vwI/AKs8GCtUk3m8xUkw
Cn9/ghKXu1eMqOwdjPnLQ8ghU8yLgs8bJkg9SxAaPZi9J5lRNMBwOzUej7FSq43nvns5dvwA4s4U
bWyTV3GwdULrCXAhM7H+1ykx4jdRBqAX6IMmy5WNM4tyk3sJXLwrz3FeGj4IeAuPhiIok45Uenqo
dN4F5eGAP3vRO/Si8skeFhLZX2YOptnem/ix3FAo+5YAtJmQSR1yblV4T/yJpbONc2Fn6/brJhby
BN7aXk6JFo7npM8zgRUZZJ17Kc+5UFA2uISe0q+zBCb66IDXfFtjg6DCGTUAURNVw461XIXRV3rZ
H5IId0AA1T9CWaBTwlydwGZKa/+bkB8iaOtu2BO1DJk+dwD7UGvye2vSIBEJJ8Zvj8WMlGDiEVxa
ku+lUK1TNQXb/1Puts27ObQXjpKvAxkVXF1aTxdPO8vWqLSsHO4KOLxS0nOi+gkkQn6ltGpSBpSv
rQGLVt5OVSrTFAIkQ3Dy48LjrMCIxD5FRGjQFoO/qWZ8a1JK9cRs3a11eGpS1Hcl6fzYZHyjtcGt
j78XHCE2WHg8n05fwsT3l6zu90X6/38CcDLHAI8ErW+WK+YBYZ4BifXdELOxMc+2mVScP6sJ1dSJ
2FWYVu4hRraY+gc4Pd8Rm7Qvn5y6L+Mk7v1LnGggmLHZOkfZySXLTeZj3htZJmmamnmKFDpwnBTf
f4SdqVka6A1zKPsjyui/eN0agw+92NdJ2Pxkd/8NZI/3UKw6zAdzWbu37uWLCWe9zYSojjWz/SJB
Qh9Nm9M7DKbXiu1SFOgC1CvZ+vc01LZk3KixTIG6riVIfH4qsd5xO5AsyrySvq5nP6wUM9T5LtyT
APU1oGJs6V6hpqCOmDOX1UfmxSF7POIO5LVkAW7Xeb2i9JF+QNvbk7+CR0UdJJBiRrE2GueYo4U6
ZbpY800U3EcfM44QlsFBbq8w7Cr6ZchE/YZTv/0eSg87iLWThqqby+dNPikXNt/pAanfjbQRY1/I
ZNRIQu4+b6wZDrT0MB7X5RsonD0mwb8DkQhVi2EiIP6Pd6i1JORBH8kNx+DWbfUviJYKOoEd4FVJ
nScbEfMP0jK47FJs9Xh6sYTnBrwf8HBFJ2V+avSItGeAYORUVGcGGhvOZuMHecLrKBhgYKpcMpQs
As4IHToIPM1fMW0HQLeMpvX8pI2eL9pLdRhDORJWde+eIJRyJfH5olzdNI/lNBQMY8lQAmGioln9
Qb5k/QOlI8JCVpwIyxULFI8xCceu6/E/KhxLQ32IfOQxfXdf2SQ7IzTrNceKg088d+e3vwdRboH6
quagVQfhmbRqkvsOrIKyN8Uu6RqIF5EAfZImY3r5eApWQmU4cjSAvQzO8xsr/3Fw2hx2a9+NHtaX
ZIzjGmtPjawEZB/iRlnj78cxGM0Ct95A63E7P4Y0+vVtAydQO2FJ98ejcig+SX4F1a0/y6fXoSaM
BVpLeYgS29VHw2tsPbqD0nQzPzQ78j5eid7+KMC4AS5/mR+hgGhNUNar28bgjJhid/gVGUrfHWo6
H7TX6CDf90jbZBb7P2dUYLT/Fh7cGieldzhLIx9c8iad4QNVevFKS0etcf42YvgOEWqkHheNnQq3
WAyC7Mdj82wmKmO3ZGWBT/tCciIvdFdRHmRyFOGGQ6qsUWFhxngmTQBVUa3xZ74Bu3a+TJSj/BUT
AX4PsRjZ2uwTsfD/qIZkkfpNa0Bz3yV5aaA83l+gL1hsjO8G4rXTM4wSz4DsR8WNG67CEQ1avUpC
8mVsfLY5b1Wwt/tGp9o2JlFCIRg7P1OOZezxCOVKaBXVc/cuokF/x4igklt7zusV9E2V+J2fPJc2
GajP78wpv2sRFbZMvMPzboQUgyncLzzpTob1EF1QR+uvhKa4V/JL2Bk0DQB2jI8rYbqETnrHsGck
WUZL9npB5ysGx/IyAcF64p3ox/lHi941k6NdZzLa7cSNPREaNEFUlcETWHeaJqxLLQCZ5ZApBE51
ndOOkEnsXG5O20LRK6i8m52YG2W7545m4OqCRRpT/KMZWPB5P3IkT6sJfbz4oQi3RcfpAIjGy5dj
vrpxlFexZY1YMUCiJUfaGdPbDH8gJ/G/ER7QLiTnldgpjUwE79gcw9tdDZ6f1oAWxvOiuIn3iFTg
cyBInSsUNH1kbqrizVzIyPZqFU1K+IIk+n0po3cLfs7CsOQnbRN/rVfX4O6pXPNlnci9O5KOBa5k
vut9VQewv7tORR6lzwNi40bNkDeuHSvzsk/q5Ha3Tvtsr/QVKQEodTvkyWlTnRrf5U9s51gn37ne
A397nAu90gCu2vB2Bu0bRuUkSaFQyj22iPy5tDFbDkwdU3lw30How18F4nqjE6fWwWH2tdiqFJqY
xPbDRGtGhx9AtivXHhLaDVnu9BkET+rTp9y+THrAQI39nEgHMneLpMODx3DLanA+SIcyPLAmkoi8
pabF9SVxGa6kkrC+MLnoUmbyI3zk80EePAPr3y2o2N7TdxBj6/6uAt+Frd4HygqdcPlIee1zrxQM
ps02uSDT3AF/5Jh0AgGjrOJPhl6o25I4JPlJBmKobB490AspBl/3fDSZXp6eljfJPs6ML8pcBooN
5agWs+qluvW8xSQ62Gjp3hpfTKRtYseWZfFYeonD8WkRoQ3qPBWMyjn0tXFEWIs/j1pmZWu50/qu
DObglvMrmhcfp6bu2hDAtFCjBIETA2CSu5YvIHKJv/81jb3c++844kIUSKQv/kE8L5rs8NLgU2WA
ps3JiRpVAbZRdF2My7ah9VL33xZ01i4wH2GaacMXsGu0foW/q+IGh8zLoR1Dkbmwy8djsvE4M4zE
yirBUPa/hElP5ovd1ahDjVUZLTW6D2dj6TRQpI3jXDFW0TpUaw90EevCBowy7MpVb6TENHHzcMge
U93yVZkJ5HPev09siokgfLcQ/UxdQN0h7lz5YeBOwvavJcGnVqF97Wd+ZnJ0/T5CthF6koAvRPiw
x+v2/ewPajLRuUJcI5SDWoDNQz+drNbtYrzgVH1zPxErzkV3bX6cEAdrMGYdvj2YUPueQ7nzVlAM
wRvrfs7jjSwkUQseAqf1jO5tCaM3bzvHMqAmGudnleE97hAXMFaBjLf4VsIdF3ErIAENnbDFu7Wc
xDLN7QQNEvtopN8Dosgwb6iXiYqvgFqJXzORzsTFi9fxPrrkW9jSACb3qwT2r33Jzj3YXY0XCBD0
K+wSpDL8DKarbdoWWKO+lg02pfeLg/JsYx992hkRC1wh7jr7gCoVxwc1pxcjbK6T6PIEIhS++SMS
VBVRVkKSeuTNDoqlIsp6IqXES9fiGMXZz8oZ3XnHLqJffm0U1FdXeGdps83qDP/dCCObfhOIM4Yg
Wy8trpWCTGchc6J1+hS5BGEuyK4YbU6Nx42HC9uSbRzKZjpl1UXThpH927JIP+zjn6uxSzoafg+V
JxfQLypKZ8Wzml5+Qe0UkrKfyFsogijtEd9TA5pT6Ie9FO6QNjZzn44P9kPo25ynSQK60CoIDCYC
Zk/oHW4G2NzuH7TQBaF48zTf7jsDP6mxEKD3d+ZVKtAaihgThP8YsGSuVzs5UVJQ2R9Zwu9AkEfS
cp/2l/Vka+0//dAhmdiguPXh1V7ZV/GWQizXP7UiUBonA2GA52Cv7tXGSnRihhvW03yQXV94Yj14
TJ2dNAJtIPHlx7gFhq7AYlcYGagfCiL3OWML+WMLYKrTtL1/oCrQ62oAtO7R5JHEX78WXSJoLQQQ
vLe+E3S7jojfB57QbLqSr50fXeISXStgNtupzTugq80CpH/Mxw3Rdnu+8c9EmO/hVDGDEJ2dyiDZ
853mIDHtGMYV9YIOIh2AADgbTqEu8kd9pTNTiEPUaWMoXRqqT57PobnkHI/rl5YoAXM6hyZrYoij
4I4tPlDrsc+OdfO6idk10L5EN+hWpneu6KyYg7Kl5nLIUZpVAdFgxoJmmi6O9gwwCRSQkxlcae9v
z9OuJmFf7b+54zKiq6w/a2IORzUOegmttKFnNDQpOTI5a5KjL4CmsnZ+MRVWdvp5HdPFDnCO/2R6
eOU24G7gNf4SLGBNx8bXjplyVi4KQ/GEbyqkzOcrlSavf3NAfsl3LROONbQSE7xbrHOtilCfqFPY
LlGWCzu5eS7Uiyzv5fckZwartcVGIMfRo9TUlapzsm9kxt9aT7G4rBAXGSk8pH5x65C+YWU5YdbN
2QlRH4Zx333o5QjJOa/7nzKshp2ig7SYlgm40TiwPjdZbdolxGsf+oWQi6ZiXekssZxPYNd2LV7x
41G8q7yuf/JEr4jkgf+h/XgNUii0XiY0BhrDvns7/fcRMa8LKporEiJOTHK/mI222BC12sXdvuOm
Qgr/ahGpjNZPOxmxrkCre0jgqDtn7+ZYbWoFC/+VDwEkdo511Ukl1fiNFPOdoBnsaCnf+DaVDaii
YMmW+poC1IcS6VmadglO2yR5mgyZLgloGY+CqskC9ADO77OeVOKs/nAQfYvLoGE2WgPKUmo2f979
yT428OEgRoTBueXLJM2Edh3bni+c/5JGka0Ua97nh9/Q9yMffcnhKFN/pfUFKE8yhBi+HMjwJmGI
w3ZlNCYaOUQc/31PFvuOu2NuFkHl8naWULn8PH7kgwvgOtlvrI1a5/Wis5mBnrHNu/y5Kbw941qH
l6U6WXC2I/woWMBj7Gqo732DN/UUO32jMmkrpnGFU0DIsdLMRwz9Xjt86RAHvp6Qx74g7bbOxLrR
d5ceMWGPPpFFlZgpPqHQECl3Tf0jeTPk1+jHbjXWkegvL83inaK05rNhhQRfaXTKCxVqfMUwYZ/D
9Q85iiciySQJx6uhM8yBe7VmnfFQv1pczdVwteLZkLtR2ahYWWX7rCCld5vOOUxn2yAeDp/Anar0
OlvCIpOwynd127RleXWOJCIolRbFX8wIXfoIa7Qf2NfDyQu5WDhRegikzpBzKW5raCCWG2uvoxDg
mVgfkmzC+oWf223UDK+R9xB8yEvNB3v9rvrAeJTk56wW8Z1pwTQH87q8UmYhvljNlMMRrvHaiXum
i0Cz/9WT9NdSX/xPulmB35HhkLfCZVkqB3Rpe+dDiQ/dbroqdFlpXbkFAHCzXhEtKXNicwQmcX5G
T8R+xy9+jme+B+u9RN6lZiI+c4sV+vJcr0YgWrAsObflbH76Z4eV9P1jlke9vtUGaMmZzCgLxD2i
Xn4dpHsfeFVPjjuogziEKh5bSmWjwVX4dhRsaBMAEcySu+m9x43Wi3nIHzkcqYcypW3pQsjJBBmm
Aw8W/V0SVedQQLB+21duwITyq29Gki2JAKNkAq68ay/RhrEqASjMGAJjej6Q3xIv6eTNfmg6+b2U
NVoryPj8tmFM+TVU+pKg3Jvka0HjiMRG9e5tNPEBvYQDhshnyyF9ArVWKs8Q/wzyjllbG4semqW4
3L1beRzYj5+8jQCaUhuIdr+U/3FWrBJXNZah30MxHwVrkQkDpHKQbuu5xHNaIJrwOQJo7lRPF+m/
z3YL1nR/JaTMEPvoZ7+5iIgFm+mj9AeGyYYe7vhztzS/dnGtR5wrrVmguJzO57y1pzDn/Az6lM2N
pbXqRBvZI9RkpVLXHkLcOnVWwhQnMEbBZxY2UZw3eHFXhpbIM8qcRBF6cp0Q7zJLhkgYlYGj4Gw3
1GJwF0sxlXHn7EEJ+Zgg99ScfSjhQXfNoQkUdvBkDf3gtvMYxZoYv1zoqzO6HONRi1+g73nIyciR
HEI24meUx/putN9T1a/zFDtx5uXgw4pS2nHrTL6hkev3S0NvYDJn24NfFNbj+BZO9O7rC+618ExF
rbHrf8x+6AlFX0La3WIFOeDLYAvhEeSyk55EH7JrELd7+4MXdR3ldwXbM5bZxmOB7xNN5F+99wV3
Erft0F+P/PGQ7+8Ui2nfTHs3pBpml8iOAWSDPhXybpra6Nau4HosBUBArD1TyTd6ahOPVAWT/esM
9EsltFTEzRTJMcH+kDYqGkdMXOvaCmpuCs2YZlKbnModwg+dwQSvh80o9T0AoIfJsoG0MXRUV4mI
2dnMP40MaB3aDv0OeH+pyruv+2gY9mHnTf60oycCM1CDAu5pY1PR2KrJET+LPCnv0v2+q0BxbqYX
5ilEdK9T4j+YuqWMEcIFqx4v2J0gcFXgm8a/rolfR1zQ5OXzlp3zLTgzzGZc7azK1+4zdWW3VWK5
rIFN9BGVZbiLiKB0iVWto+Ii7lvuYeWd3o/GjjL/XYfk7jPvqeMmW2YNIqg1ck67vBXXwDtEJ6Ig
fYsDSAp6vuqp6zp91ZUdtbI/47KPKWa8oBp9X9qfXcNex2KSk8UYNJX3bsMuBqzZ26CrwUfPp1Mq
42BNuoFEAelF9mzI6Fdyy/7rqlwpvaWWmEBBKDxS/TysRpOYPEdp7ed1xUEC8/zpUZN8YLhxgOxg
g5y8HiElqpnvLXT7iqAJJnYu0uNBzNkXXA4fzFLYEg0Sa+IGJr8Dv6DTQ98m8DFcsoxiHA44Bb8M
QdNMrhWOgmtqwHLbalTGED+1trmFi/xMMoZs6fdLEMihfYEe+aVa7j/rFb1TmstTKXWiN0h/I9m1
Pp3B6DRuXa5DXn8eDI2X1+RA6YvUznrtiZliHWka/c2+I9sEyoz4QFZiyfGOugGMsE9P1fmwmHWr
ncnQFxYfkBnEYIDUw5ja/32Ka3yP8kz88oirCT3y3Fx0cBOUayYEAHi0/mSTeHCRE/hx6R6A69sn
HTDF60uMDnGNZqeZiHwuZaBRsocGeahqLXglx/vC29ACzbzLrc65HiKySveQEGdHc7M8EWVS52Ta
YcFuuj6Ibsg1MM7N/JvFoC583z+QCBn7jQn0ojczCYv14gBMbcdKrir5y82HIyhIssVbA4e+Ze8C
tmqSFTvABIR1p8jBDJfMagFHQZrfWSGV1zW9MZKeNLoswvOUIR1MTKjZ94Wd05RWfpH0ueXUIxkQ
PtKxF5yUt4DKukofLvhLE+FgSXCxM0c5VKnc8zrDEU2VXu9D/uintKMfylisHgz+uuIOXtHHwrGv
GizLZpNoIxynMjqWU7SOGqkohOMu4NAOFgYgAJhwqUCOwaGU/CFM1jRF3pqV6CChrHmeIkxrq12c
PzBm1aBnCR6tgOAuFsa5Qb6pD4oGd1sN0b61q4yK4w0CDIgHXx540cV14cBjK50N6XKcAHdochOX
qWl7uBKSW3TGK8MmB6Qs2CskkSdYvhrQfxIbPbvT3GiKXOLh6EewPL/2oVbNjB/zCSBeGP8rswRu
j6HYRVN32E/pvHgeixYIPJ13LETzgktSm32Bpzc6OnNlLWZQqsjI4a8j1GDHtmYLrVT5ULtoN8Ry
1dkRy4b/9SGymRaYnmX5LfRZJpppCPwRE1njo1N34IpDB5ZVpcZIIQ6xpu6mm8EscP3IvBX0P0+n
8AT0L3/fyqVHd3l5U29uceIvOp7AZm73FsUq/jxHFKp64Lp1l9D+Sr6T2UXgoiMLSjfC92zn/Ahi
X8xI454Mgg3IsuEnJbMDlgOW+XaHe5mFOVC5t4A7PHK+AZ4ALtsvVT5cyUWX5Gm7Tb4YoMOx2nT0
UwVpHRedj4+Hs1MKE0wAW2rMs6DbUGuUCBkEDpLav+hfIhvo7Sg3qW79Tsgey1YIhQhi+f3LP3O4
XMIltGGCUQOtgYTL7pgoLeMS3b4LC+LvWnrgJEKovQOroqaqxd7HTmCnp+aO+Cv1PJLowDm6P1Ea
O+HQpIqUPh+1QZLI6RgxLqINdpA5GZ7G5OG1N1HkaHGJDXkJa0ndEIX9J5cPicaoIslFxBAYOY0M
a9X7/7z5ybvVkZ2eX8+SRwz4h9P1WdnT9bT7QLe2p84TyjSP4gOJ5HU4tea2HlRkdObWW2d56Nbc
5vxiJd//4fJejSxSBk3syy7iGGocBT7tRBGNlCfD4UHYbNZsSCvzh2ZONLyv1VGx1jC+F8zigZFz
UUPXd3xE1ZrUGizqZnDgT/eR/fLbC8R87hVBHVvkHDP4zPwuGrTClJCNGIHlnN1CUkuBA1tdlX90
FwrdtDejAt9GoOC60UPXV7lq1ECpxYJSWFWIwlQ/KYMAtdY/4O0RClegy5OMNSfLbSjw4VSknC6r
KdheLvsxu4ss3fWVtsCMA3FUHgZnX3a4OnFayQAx5mpN6vVkjhEDsvSMkDdbQROFjKGEtx1wY0/2
cLp37WIuN5b/Q5cCmblchwadA1s0kShlZamceBPpSYkWGwShT6uJBGNlOlPTabHb+wEtZBlu+B2W
UaJSXA5ibfrXKDhCJuUSoSfV1Z/Dezc49Mv+4rOd3vrSYUInB8lHl85VDRSCkAPMFPAsShaHEbPS
uUU87acsAGAXvFPOP9mjSj/th5pYFKSAnkfQfXPM1p4iGIkjkGLz9ssa1C9w0CBMYX/rUCJRLUKj
ptH0yJ/e1INFDIyJUMKDpG99LYJg9rojIJToXKU2K+HjmDp7SfRGIWl8TY0dvPOfeEFm60xAdq2j
pLb3iP+vMpWuQjFmnxQbjC+zKMl5sqISEhYhKdRYpHVOKOL3VPv+PdmK2D7PiMZwH1zotaToHYsz
rn8WwvQBVKYBWmF44jfHzmTTOpwUqZ3UH2u0ZnEZFh/8pc3juZ9/O0ssl6P77diARi44/VwKeK/L
NKow+pzjVavJz/HZqf58ztaHoYxkPc1xt7GlG26Tiu2hutpVkBH7kQqxuHZ8W3tUj8tF2ZE/QWVJ
sc5p15AKO5F/LVoCkDys1/pAwCieS9fMjCtUUrlJhJ8cttY0rklQBpV78K+C3b+YqMRc/3w+T0E0
92z7t6On/CqP5wlQ7o382G5sZYvxitng26uIL5RTGqLPB/b6b0aTxtIXhzkBlxDF7CQxF9lgxL2C
KuT4fxPTaq5yqrPeqk4wEK65T2HlYVoAUK0MyA9a85d6rAwtZMPKREbvZq7dJTRyFHfrufT095Lz
QXLP70/sNADQKVeeldUFM+C0Bbc6vHPZXqq+vVvcwPBIyFwXK0i4slqUrVxoULh5nGzIgIAxYU3F
dIyRVPkyBJLLl3DX+7OYHo6VqZXXR+8HH3vRospycvc6y9MEsNl8/SI+IZaTd2yhmJ/nsXTAtC+N
7xFWxa9hEhzvaePyOCaS8t1006a/7Wfg6w1gR4HtEkN3nz04jgR4M5TDIvoEtA5ZIoIPAiOAHBX8
qe5/ZofkPRs1WKtMZzUy/zALDSsooEucxXCmmhlDXHj+l+z4Dzmocv8LEJOwraJOMyDlIJMX+1av
vDHwOkuZbD0uO+TjxAOUPyRfm6v3uoBG5w8Rfwdi1kNRN1lMVypVjGgoCeu0VdI4xADL12Iq/0CR
ouU60CWLnQzErkeJysJgx5p7dPNSZMxCcJM3yy2SakurJmpZwXfJEJIbc/YQEmFmtB+I20RBkRSv
OVW1JB5qdj4CtxqN3J0W21A1cs7eCFi19XvnwADlmIEke0dEyubWZcefqY1OoYYWfcSB/UernBKe
UqG5GYX2Z/Tx2Y0bvVU2CMAYl9oAULQ4fv6pWXAh1XODjDi+ULfIhLcCOt9cPKPA5il09HfIjmNX
XA4jIzgzKutxjnSg0KYMmi9/wsxyA4v2VwbR3zybUS1c35cKH9cVcxslx2SM20DdORQ91UmDm6p2
BbXo6Vwa7QV1B31A90uVWPydepxlqYAqiIDVhT819KnSEvdN4ctI/Ccydw7kqPtAHlPlesHkKuJD
IjdnJCkUq9gEtVyNvN4U6GQFsvmmj70uJqR1FkDU+LDLFebf0EiQdhNqZmzBAoDk1Oz+DOTxBZEa
e1UuLV3+vEydXVJdCpu4E7NwOltXFBlwYgmsgtDhapSjRuQ1HpzmLdHNsB/m01uG72Pzf8WNlB0p
fxyFkV4tgYhVQ9mEoCXCimBKiXBZnAKtrTDd4HmhznMWgoX4rJ45THdTqtzoYR1eLC7a5zLOfq4r
A2El6tXLGSmdBxPAfYLK6LgtAp14KRHKSSXKGjs6dkKvm9i1GnvcCeiWhUNswJYkn143HMGQvvfB
E4XPZfvG4aet3NoS48RCdhANFIHSvVapVqce27wyNd6apkr0p9/Poce5QFALcC619Cs/8ElcJAwO
v56F/fOwQHqchLtVwOdtyts31Y3k54Gv9xbJ7x4bdpM9Ci2BP/DEu0AjrO1cr/4XEV1lwmtKfiwZ
SNpqk+RlyZvPDuD53mwyPHHFsKTqKLLwJYLvetaRHH7Nl0tr2s17MCHAAG+msRE67gZRplDpbmgx
Omz4htyB8uV0QzSCH6JXR5HlPD/8vKejYTtqhyy/szX3Bx7Fk82vhcF5B7X3NSEKeiy0qEL421bg
d+j209eBr38ZTjnXtQMPsSpfoVFZowDkrNltk97G3x+uYY0TIyo7cfRrMVfYBuFCs33fxdvk/gpg
KVdgFxhJ0nWU7Mt3Pwd0HirsUg6f0WedtbiFf03WCh7hT4TIJE00rHn1qTF/Z2Q8kfxVvYViFFtc
fYc2rKQH+BjAHKjTWsRGX/ujF3ATGBh5l4VcWGyM+1R2sC65lsGOSo33I8EzUgQa8DwCHCIrGj9n
aHcZOuDS/6uvXX3o5rkCSOAl6PTXExKQx++jg+91TRZ70mdraez7eBaI65HwJsu1Asjk9QXpIVuZ
LVaVh8RMwpDq68awOiQI2zayBeuRYuvYzKgk5OCC6uaWA6hKQpWcmvKoulLtpMCnr2QpIdguxdgz
ivmS6MzzMuCTBPGeHfAgftmwmykR4uqVbJ653/BacsYP0CroTsnT/vKI36Qp9dQXASFRv05WBUVY
iu89p9bTqi4kdSUlsACa9lNX5AufLlJ4udJpLJVC8q5UMysxFP6VGkWrcj9hHwWnTF6dm9gePOQn
zbfgxEwnc2yZU9QWqKMn4ffEqSNe4ogrRurmRm6JogQxdhKj5bbV+5xu0vIb/LJ0rChFEzH9rYoJ
vjGZBnUU5nR+0Xwqod1mc8RhqfLjqZgsWAZlJlUFtkA0x5dAovvTpqw92rIJskY42K2qZPvMGRvw
Hc9YUhqQwhwHPdgo3Yat9kINH6oQYxTheMrclcaF7oZiQ5JZZHzhMF8Nf56Du9kbpUdf3GydXOCy
TxTayYmP0m8jA0CpTj4d594Wn/sbLHlWFaUWPIwfOwehgeUiVIY/4f8vM4VETuzpZ9n65YUWEopW
xDbTyWKrkoW6UYXJ/QrqVw3JhaS3tJ/pyi6BO4OY2QYbG480aD+hYnatZXNAjcuwdQizpoL/Yccd
O28g8ksaDabd1c5FlzcAj6ry0MuYTDBuxbm6cCbZJ8I+2vxxSJGTRJ31PtnIv1JuheQjzNmwt0mC
hNXwac+4oDSApyldpzN0N8o8TXp+YL4Xw3CSV9NUOZoIKyne9YbwdKNjNXToSGgRnLHr2HqbClGE
7Ksq4SmDbnYGRvg1gaiW+wuV9iKE7LKoZ0xGDikfpIdHRIWvAJFA8OpA1o9XbdICMYKwbGx7WXeO
BSVY/Rd24VZMqFkkJNpZU6iP4wVOk+Hp2XeoCvukAamwYxeuBuhdBum7ZeVy9Slie2m6MyerLxbu
6lK1n3njh5QPW2+Vlgq/b55S24MVZfLSeR9/epHSIsY2pkcw3K4wABFQB0ku3unC3KLv+cRrL3Mr
aQDrLFaGjU7aujdWFYgydR6yS8/kYyeZasL0Xfu7KEmlHRFLFJx3w8cGGSN7+gv55sHzXTsLY0Cc
CsvNKPaDy37p2Ll3ifCPxXfNULXMbi/cPzy5CgIf98pbko4RMC9A0/p4lUFrnMeME/VZCXHyeIJD
Jg8wDLuJfLfpipMfUZJkcKjWUYV+GHy8kbxpTlGLa20H0r5flRcttoreYMyEc5z5XD2I7nybROki
Vz3cxgTncEI7i+XIx6yZr2Pfjzjx5pYQhMPsve7Dxaxuw/1KCBXwPJ+/gI4wqn0b1uJ5tg4D5zMB
0onzlNQULmLZg5P9hVCv5/WnAqSmbpWXxeMsPBerEpbppr4vc/akbtveUQ4VoB1WHdIGJJDJXGOL
AS0s/opNYaMskFX0cBLd2t7HWy+M2yup7tFQARi2pltGvQA7+hrSUBnRR6Qh1E31F5f63IPj98/f
4jj1OlOcK/6gfmxbu7c0WQgE6mJRgQtYcO2X3vqjx5jW6XQSxIO3Nc84n3YLR5oaRiwJnr4JTyCo
JktjnVU6QglbJAyaaKD0wlCWcINSGOnfLL7L5MZC47SYW0MS7MAwNUFLto+Rq/VAsiemWCGF8sEb
NFJGqcWhANtv7892DbTNHDUoc4/639nbXe3gMDJMWhhmzVceH2Eu/pfLFoWW1I7X9MREQJMLsB0L
UQ4gq4ft9kjsSNRDJxb1gl3KsO6if9grkOWEiE8qlauqjwzI3krMm57VmOW4Mb/hmTDIplrHjciw
PzycEXvyuo8ufYHFbVE+cQBE5+g9yCb6eqADQQczCkFx/bVKiuHlTMAaBjod2/gctNkdmpeQYvAj
v7jPGLrDWFbUN1wXKiMUcPXFIXyYQUxZ5holPgBXnJYGj5p7j4boZzogW/h1pPivPq5NBj2dsZz3
n8T7+BKj1I8t2cYO5tZCFZIkFXOaXXKjATohRww2QAlZrBuAw9MTl0iPlS+/74lZGctHii8bpJtQ
dcF+RxWPkkl+QuVAVo/TKdEf2C+iAg45lss7mVBjtE/aBfH8TXcmQdkwLejBmv1cYgkY9YxUXTA3
X50PM1UAB0hKQAPiRM0TgxxGNinrQSeK0XXD9Nv98FiGABnwe+KrXUnkGL+fYZgr9r/BhnxMPGMa
QmOr88umbOhL6E62B4eoD07BQKYHTnMUtra+FY/tFhzIuOhE1WxR16oJtWs3mJFqCStgO62n4nom
0l4b9j/FN5xeY+TQVzkcyWAnWiqu7VK33utpWuJVXbkCZRIL8BGG4TFVVkTiD/75XPf7BchGtnv/
o0PrZOUI6Xwlw4KUfVMGqUtGdhbjShqmw/6mjthc+3uBIKp5asO3dZBHGkRdwDD2EaBm1524aqqf
tuB4FEZXFMzZ919+ZUfXIP5kQkl1zynl3RehK1ov0m1sCogyzp+U19IFICtI9ShlN5iGICbCBr/S
Pqe/1zjWMBBj3OqL/5zSUlNzWDMT534fgxqrVuKGQRypORuwYYJ4Fwyq7qfjTq14VSsVXWI0MDrs
2fK0suFHJG+1y7SK+wnph7cChh4KBLFRQR/Thi9IDl/9/JL96cQAgshgS1arcLY8XNn146QFkC1n
Ui90r4djcLigb9QjbL/OPeJiB3ATMRRoOw1+6wbZF9m23dKhOxZsCg4bwKaJ2TMCuzPTQkfrmdbD
yV0R77YrJwwMSmNeHH4GV+mzHTgr7endr5X9pNfYlDmXxW10GLqjOtQak4Cyz3XfzobpJ+2NK3PD
6ZnNmfjaSBqyQvMFzoQ5xvBoWi3bc/5jErV3/JXf1Y38pBSrrqIuCXBnye5SWxTYGpY7H53PuEae
eU/V3JAksvo4nzTQz2YFtK/DfoBDb5oRLXdXBz2lhDuo1b9Iqa396vOJm2QsY3JfwPKoC43KIZG3
TE1W8qE/NtfN3DM1m8dO/ktQ1RZ48XtEh9t8F+oS2kpCCafFLugpm9gOJw7EJhWf1dfZ6QoSa/bE
U6O0SX4cqlnCx/1iv7XzpEGXStrMiME8MaSVcyE466lO9QrewWMN3Nd3+H0QuxLGoqrmyi4piR/d
XJEV9ly9BhbeRjPN3Ncd0volWX7y5RaMHze2clXRLwdXonomEEQWz9BeCpduYPiwddw8pYNpYXJ5
ma4JZ01SusAbMlFOqvCjcYoz5R1/TVyM+Pz3JouADZcw6+5WdYi8dM1GyXAUEE6aoSTnXrVJvyxs
tj9M1Zu36IP6wGE7+sLhztaotuypDyxzZmRlbzaoCds0Rer7KnFKqMJOUVsLn/yMyAdHNAFm0Nzp
toGLnwUcsclsb6RuBNXf1cuH15Dy4FgBAWIS0pohZg0oX20+eA1aFnva940Bmaw6aMSvjYWb4vpF
6oxDOXWyfe5pHrHtIgNM5YBmTBbv+oPayKgcGd/CILVCXoFE+qcZCCgQR33lYGV/0NBiYOAVFKOy
jQnr8oV2Vjn7ysxmMCf9jsamXo5wRT9EAMF9qWuZA7xnta7M8fudGQu9Ma1M/0/KJysz0yVWEzVu
TjnQ6p/f5YgiZHd7TA48zC8+Dm0giRVo/s+4wEbZ9NEF8NDacEzqdmvCz+nOMiy5o919MiYvwpD5
dfptsmphKcxqq0OLuEYxA8oaLhK4n9LIfWpEIxBl3GLO9U+ukRUBLyWN+p/N4XFjkcsb0+S5gz9m
PRW4YHOhi/J48EZQkQHu7PwgyRgdC3GBCBFHYMsCs11P1+C0NvNzgHNtxhHIpkoi1spOou/97utp
yvDHxpj6rByQs0Gr7pxKykc9pcWC/YbRQr0bMgKi14deup4rw0Cvgc465Hm3+Xg5gcb8oFqzahJI
dnx1qfAs4jTVjh14UE6g68rZXUaA2C2MwAweCBlMOFjQotgtBtY2R7Tb48ojKWIHw6DxJ63GPZqX
Z3LYrWCygF9TEwPJGB080VnwmiU8MqSIgBGJMNRhE+uQJaKsk3rX9hYSYUqBf72qOrLuuXLuNzHo
iEKpNvd64p1rbb9iHDkonR7mnCXzdKOJFR7FtAkOaouEGA55PAWZpYF6Y7xuDWpDhNwEzEB72FW1
E0BwMovox/BRC9GYa3l+cALN7jnW41pKYoDHHiFtvGUMKyCXUKxtfqDB50EaYF2Evq3I9SXebP+i
XttXw7tb8+8jDaUTBf17q2+x8C/TriD+F6QDrkNJeCvuAHsglejGzWH497++9e7kcXkQhMiW+wFX
aKYxtKaL95VXDW/ebgo8oeEEb4PKavrL4gtvD3bLbp4nGMpL/xjIEWMSQ1SdWElrBTGyaXk+aqJE
aPEbHkzjXiMFAaYjolVtpCWZyicBUtC4d6LI+9vkW+zBFwQZImiP1x3/5UzptevEu58zdphb+CLd
vRPgLAg4pUOeT2As9ckeVJEAL6UDTzDHK4a+XLbfU7Z1haNeGfjxukqRbX/ntzVrF+5dGUgU7cz9
uSaUQDzx9jccZtUKuBcgZoM+XEwlOOnH45mYQsTgzJGCWelbncyLPzuMa+zHr4vMjhAEckOLqk8y
MLXwacIji20/bo8bUhAdXbD1/ea7oHNG2AOKo6+OHhLAnBOrYqtJx0aIvXUfBYiSx+cUVX2TwzQO
cIuefhCeqGg4vE5RW8KdDRQmH8kCwLRN/yLbMpXi3RmzuGM2UpwmL1c7h1/8g+8HHzzkfrCqzOp/
GC4iJy3mUiFjWRKNzTk8t1Bcye+2g6ghAwiANZoEx4ItsqYcoIKBt9HewLEKKD+596MO0XldiGW+
i1cYHEjp74HGl7ntH09nKpwOlXDJzZqzeBbxh5bioGLI04/dLTC3Yhl5yZBfjs5czCSYDbO4Spge
3a+GT6RF8Cj+IBQt3NVeOUzhl7YYpuIZ0U/r7wMIDHYYbaNaXp7QgoN7Df5VrfEOK+QhK8/Nr9by
uqJHQCv2aLFKy/F4v3g/er+EDK6oFVPMExXJ383NMY3mzCBPSXZTiBgauNboxnQzE9w4sSoKNwsp
nYK0E2o4QlA6+5kqcBGdzzRAG43htcXUqNeE9/Uegz3LhymWxtZxvjumSCM3TzivWFIJ8lsXa3FU
+Bc6MsmHmKz52GoU8hpw7QZ/svO9Fp6fIcRUC394P4ji9qP9goLhpnX05jAVJJ6wzLyyNvaamFWO
A/iUwQTGLULZnP9mlIanDIzsvx7fq2U8qib7vz+8bhO6SjvDDhyXdm/Tp7WPYtR5eN3WApzHvoLF
cAm4ZVUfHW2nLdAZRcgOX1UooB+q1yO39NJMyiE3DohJnaRaoblHH4LcSPoyMIw4JvEjPDCrF2wi
WLjEE6mxx6i9ed7Lr5VZ0KKoWQBp6/9vZiGj4jyC3WL2UEFhgNfqxMWXQZ03QXk2UEH8dcXEjQZi
p8Dd0rSYoInrCLc4GntNz44N1eS6HutVctAXo5+TlkIO2nLAjK72AC1n/e09bYeWbSChrm0C4HMw
NmUWRF4yesvo92d1RnxJBbxj7iNg/R8RBV8SSERfb5/ERSDuMHaHElceUyR9CP+dohIgkUNSd7Ev
mnVGNEBWsSN7rN00Ewx4vfuqdfwYMBKJS4qfCYCdAudHWVbK3T1pa5koSOAg2c/Gd9AEdPXtr1VL
jXn5op3t1Iqjgos8FEdfZX0piJdvE+qgvBuo0tU9ij0UO2YI2P/vnn+jl9hShmMgPkNd+iamvju+
B8h1ioZdWJF+TRuY/U+/LF8cdJBsom3IpTMSm6sa/Mktt/WI5k3MvMMvfut89Ts5npt0kq3+E26/
QruDpZMiBXEvkIMPMoLnA+izvdyvAEtZei3gq34DcJ19ef6ZL7P5TpA/pGde5Wg6XXKLi91jnbdS
zSUpKhyU7d82RX9grznrN9SZbCM49ZQUzeq3GcWYbzJNwwRsbuYNIXK7p0FPQerH7TleYsqLth2k
aOGkfk4jRR6mJVF4nA14/e8LpH82f09DXHI91mbI2npzPhD1GmpYLxRULdtMYuJtybzyyr0Xmt2W
lNSPudlbSD/ggdcsdFh4F5uEWH/Z40ehGBVPi4PSVgrcXLOUV79muH4yM8wpA/TnSx+bfeNOgaxT
MPKbnub7xW7kstdSwsXvswPebRR2JyFZmdXhhdrRNKVStfVJMCGgB6oOIvzngj491+t+Cd+MkD9N
h0F5yOpEj5ckwSv5+vNuF4kVuG/7n/toq5J6z82zg/nKRevr5Cxi2EU/3pAMseGTvLSghFkZKg6q
u3Mx/Nm0XYBvlrJJH88gvJimxYlzcnxfFNJpqQkqOISeAruagSRoQ27aNNYtBIGYz4i9rtzBcEsJ
DilS8U39y8bSOsmDGIV67a2mELtHv35zruCZu60BQl2Gtj9pr7pa9zbMV2dnt8RruPqaJnJsZEqy
6+YD7nrEEbbbtW0nusAJINwc7w1QjpdQBKWl6m/eRfq9iTtTpbDsnGwB/FIr7VTbARGCgXzEnn3C
aztwrIR/TN6CbpNtLxGFh3ZNjjr7WF87hciCG21O4MUQnFiJONYP3TBhTdCrhFeQMxnU+2dm1KGX
UKHqezCDfBlpWFCt7VThY5UMmpBkk9yv22JhBys7EDLjvZOkLwKQw+O6Dqivo0/eWNr3AEyDcNEU
k/GWwIGwC7TMiVLQs+rILBc0WYFUI/uw4bYRJX/kS++ay9Uhuie2d1Pbh2EmnX570tTeiGADggq1
RDj+0b0yIPCOFrkP20s0zhMHtYLwjJ/HNlL92P5n4BSk+wPJ6zPodJmZ7czBRNeDuI+KZXwiQNZP
nGcFCME8tb7e2BX4xaQY44dXMZuc3Mu8/XqY/jDWl0x+bZNXC04o+IQq5F0dAGVwMXX7UVMRxGKV
zL38Zgt8zk0J2B+q2LePZR4KbG3vsvJHJtIpcrPyCiror4MXfsTDjGPVuxNuPfePZ2oPLoSjxlwO
Jg16bmY/ziXWgeDLyxemLTApGci3YHBTcKm9iMGNLZOb4Cm596m1GFOrH5pyEyhXEM7w0eijJ+Xi
4BN+KsagjvrayP6CzzXH7MMWU4y8vAlggLY8IDFouap4oUarEb/vrg8jO3zBBg1G7Oc5Yjm2bap5
buxtc/+iChd72IPAifeAVc4rkvbiwKWhkZnRCKQ7q5j6Tu5+vfKDyoIYzyX9FDLIVp/jKPnBArJC
dD9b+hrGQb/1DKgeE5PKg1PaN0BqIJA957L9kMx82tg0qWlEl/gBjKAadnjQpA5mGO3Rd9hF+6k1
+gEDdl6eqCajz2Bvj/4DydAzZAlfHVJU69AzEn08V9kZuY/AvPC3D5eQnjGa4povfKZ/51ps2sVY
Bxg57RVxYu+5IKozV3ZEUjTGiF1moSc9sTNIIuR8jJIwq2e7L/9tugu3JXX9DZleoRr5bv1Nfu6F
mnDDbYnow8VQYdey4Wh/o5mZFKoiCfO65Za9dyI2A2QsN9ahqV8J2/uibpOjE15FwBmEM5cOjJnO
tkRMfRARQSiYjdv3oYfXyLA8Bhmbk70RDgLEu/Mj3SY7ST9u7bVOdcSww+PprWdc+E0/Ee3/q4BE
lJoQ+AEkcErQxLKVjzTGVzD32oKrCpKD2jxU2Q5tD/AVsr1hMkHpZwJXZ/+Yt7uq32pDM2AeSr6m
3ulTft5BvCJreP38pieo8glXQ9NcO3P6NVE6PKqyG7uBifHOiyYEbIRsfZSQZLT8sQCagtqTEjx+
bLSXrZjYV9KQvidPpIG+41mBuLPFOZjIMX0aOIRLOgKMIZNd9ZyHcUsC61QLw1HB/+d3iKdppVfo
tKQJcfn3WguIO4OFGUIT5RLUHLPrByNjyHjRwV6zBcy8ZXx+tRRsEFd/fBcOof4lj5U1tQhMZj7q
55yE1Dsl+Pv32l+5ZA6zT6O2MH3t0Jcl3HQ3J+JzHh0b3jeO4yDBls09EE/DQ1eEdoNr+aLYycEb
48CH6Rj+vp4478xARpRGtC4v81tMtim1KS43Dx9jK+tw2M8Hq3JJAAqkcOaXlZQRdD6/Qbuecto/
QEshXYO0I5wjiEVXpWlymRkUuGcAJkQRoxx4r6JJfGHtIpkntJd4XSAtJSbCFiHiyOXuw7lIdzj6
vZZCFWPAu7uJBdMgBWegv2Qx7ntg4fsc4N+MNvsFvP6fB+kGwZxBp3d14cCd9ID+0ITIh+tf1m0F
AhzjJ19l6Y0hIQtRV0xS6QgIy3wQG4rT6VZ5GktYxr6mLenlwJo8lybbrZa3UiGNgcNkHmFle4PZ
/0WGSNXKGgTlXXMbaHxydVvgH+r9XVlHguMAJHBUVPHfkzC+6SSRQlfxMjsl3C02T5/YRQv6zQWp
opguUzFgfG0AwywECAgXyFcDtJvXCxtYssJkDJsQD3eq69LD+v+eJgg3f1h+BBV7KwpGmqxrCORo
rzUs7Gxcug8zCIg6PjDU1NoqhKl6aeJZLRHRkfyAZkmRsJADshPQPU8ikPukVPkF2QZyZlMUKKTf
T8o85lMguL5zJlK5uK0N2MJ6leXREcz+vAJh7lH07vf3B92+U7KioVO1nyi4cA5DUl4eKx/LbEco
9pDIayWOalPZxroA6IiqYN9JyOoaWx4uBY2m+VLpEqSICZcvVlt/Eb8Ac6PbD5/89sL8t4hJZzjA
xBcJx1YgyrBy48IJoUHNRv/6ZqZEEKLxvYQgy5HwlTfAHzyawe8jlStgkiNWJczRaASR9VCEsWkH
Fz85H1zLpv65618ULyia1ERtC0lPXv5NR6oZuZXasl4xsQACuBH0AwUxHNF8nYzFwTz/sKIuehbi
K1+N3T5IYMiqDUvL5Xd/oAB0T4SL1kCIAAJPemX9ksWi6OQgwPgds0OY14NHGXwEqtj5LuqEV+fL
5SEwZpKUcnZANR2jBqsymW+rAt2G73JGiZhFfyYw9p0zoR5f70mO0aInw1dphSDsaBAoUYIdTgwc
EVCbSuD8t3d24g5M9jAI+EQzQHwsrq7qy+27NxEuI8A3yjGel+Uu1YQz+TQVpr3RwHxo97tTsGiM
JcxtINcj7CJTVTyxOCf6ajKBH31HoDx//Sg0hCtfqYk1mmBchcs+lAwzxC0SAh4JwbsH9PKnorGn
1gCXC4Z2Mi4h7tqmI6YH3cjVcG0Zf98440saojKuztqn428mNKCxi7PkMPWQPFDbFZnMlqfGtnDn
/qusFAgzPIScewyepzzvw/7fTlwE+p5cLsRf2ztwCVFhdEs5FgUrDM0qwwx2CyeJGyG5IpUdvj2P
KCyXDC1LLNsfEjBvr8CoZFTekTGjySvp2qkKSjF0R2VAJOdsHpeTICzqb+uCRcR48O9yIA7t4GAE
EtRlZn3HTyveAxpV5OPYUHOog2LN5r5VHFgDihPpkmaHqndKns3Wgf7Qki+NMxAU/xOf2lyFU5zJ
195BDyzYLL47bnsnD8o1o9f3NhxdqjJYXBLHhuToimZy/mSn3ZSBF/8NuhOVzYizuIgRyED3v27N
W6HzkZCe0rUHQ8K+NxuRh95f8aGwTb7bk/rWrbt+fD1s7RGekBs3ZeALQy4++6T5W7SftgDjtH6K
YVttwwHKUB/o8skEMVL2D41y7bKYWQ/yRrMYVYt31TSEnKIOqp/Ckv9XDhyW4FV2db1w4HNv6NYA
zThRLnstk5a7wmudwovHymo2e1pGSMXd2Ky2QXoQw2NNiJni3o0AXCErQpIWIxfsW1HvxcmuJBAu
qc5/I7vYpgKMUPHHh3/C3NP/9ptJDlxGObvp+eX0lF/+wV66O83UgOYWPD7VR1IL7w1eYYUYNtuq
qpvGGqN4fo5C7cfMxNk7OfRm5U7o/wYsQ/0SF+/TnNt0wRSOPwb2mksJT5FjtPUll/vJhtR7G05p
tDCYemY3x5KFmY5ekjcp9ME1jXSDTNtQl30rf9A5ziKEzMmjpnCYu8OIBgEoEG/JcOZy5W5GyXMW
MLZ2HPR1tYDx+O2Agp/32uHlKKmkhvpeeYiM9Dk592mssZr59Zy7lHwvb0K4YdqB7jbI/4/vYhgJ
YfTjZv3No73sTCukIdTls5vNNIHBH7FyJVjBt15EDCeVff1QC8qr1STXbuN1YpUc25oGUa2ZCyPM
V2XmQKnAlPkyoRP4WaWNAsPO3mXeSTJUnmLF/qHDSLq5L6xiIBwTAz1VeYtLklrHcQO6Bsrr1XbG
PjmGHfaeC+8Y8PAR4FtFtyHwxR9yazhfSE6SjnZCDV7DWD/N7v2tM6MimsSu/OPafNCRapO/9CNl
yFQ25YFgsatqo4ViYFLgV79dQniBQ/ESxNGtodV3TcwfAjdRSVQR3we6jTbHzWu6wwwTlsQ8E5AZ
sGLeESdHCp0/61+d6EM+gfphKnSLZFmMGe5XPBennwSepn77WXNC7zRgFiYPPf5Is9zQUS3DzaMb
nSXz3BYQOke4/vR4QBDaYFSswWbE5Bk4rd9OlsJNoL2Teym4MQ2efDN3y4v3dGaOeR4Nb3joG+u+
IwVWviBHag2JbLlSIoN98APCnzTiMpEL44MOg8XULA/lOxQsO/nDLcKfD4jrLVoOIYXmY9WPJRmw
bJMQP9gALuqxPLm2wFMYDT/KDhh4st9yU/ZZHHfW1mKYul37x00epstLKMuTbSzPCzSzxkdwS9Pv
vnpvdWZWpG3Cl/ro09YH5c3Kx85PC+cT04MePpbLpQpV3l9q2/Mk23kxE1UMPZzDICec4kxeLQvS
US6u7MlSPxB4JOY+z2HiF2u1AFp0qiVyfr8cqBu9SHvKF4SpXAQnkOmmXKZqEADc+UghPYYfbjsZ
dPYnwpaLy89YAZnB0bxdnFzsd1YdEi3TsbG0FJhOCKn1dBoKhzT2YSQdag83WDD/CZcm0SPrYfng
RtrikwwLZ9WlLzG0nHWfO/KoJcaYpnWZd3XS5SDeGUr5IAxIdPtRvVgIIMf2ZJOuEgy1Dh9/qwFy
IWrqgjeC3tut/SiuWuOgvgNwX6RIyP00bo+I49wiZpCbgpUvzx80Mfb7evET4yjMxTNhZehnaAHp
z2KOh//RT47W7JzoyiBLHpFiAuQBOb+KdQXSPCKk1KCNZKN5J9wkmFpC89ZsiG0nx1o/lXU1SKOC
maNaF2dpVeNtOLLS3FTFN0lntkkUPw3W60OM+1YntWAt9y+wS4KbI+R28A387kRkN+9jH2gCMv/K
eJa9Aw3m7/7NEuQm9FCkwGqxWL1iewCwKIwRI+xf/KzKunihuOvzG+WrA26NMhenw9ni5UY984nj
geRZ7LtpVx4zBZAwM5k/xMLKWK2+livl6f8fxOOyp0u7Nn5huPqcI9QZavr+nRdz3wuOknDUeUkO
n7fBGOkyuw+pNDPa8iqAGPS3A7vYQkC8PMLGt6+Ak7//bWZ59jbT7Q6yLv5ObYXnn/sdn2DP/6Bj
OshifJUcLFQu6N+Vn5EWyRww86F27DHQorgeAvxGtHNB7xvYl2EIeaSFuNejoWaEWLSZ5g/3wIR3
pSyyr8/IFgkdpUcuZ3tKKj5v8DNMRlHyCsUeuylV3KmUhUexpXr4q+NkjNF3lnGDTJN5ZcT60YHg
ZUvPmD53QvBQ9j5oszXtNTAvG7ASRbVIA6vi7DohUMw/Tr1wF1jPdwRtVs3iDmxKLTgjYyCeGvdT
ETNfXLpQ2smVZHy+UCg98Plj9Pdw0j1CCQy/FoFJIbW+tSMDf4ubjx8c3heFvjSNYNe7Vxu114jG
+NyBd5BBiP+/zP1yt0PMPhepWBbT2vTT+uBj81MuuVrW0YJMMTyF4xxO5FF37rqpcsQWT6lc6tdA
IHtuNvNFWOibYJDw+OlP3NM0erkh+KSONwNaGm2t4a1J40NbX0FRpYYKdJlFNKfFMWbXNPtDEzRR
i0+dHgqYHVHGV4ya0GGz7Gt4nKbDuFXhPjAxgNVViYS7H99c3EB4qQ13Jk5xHptZO4xcALlqHu4A
ZRddRdpQAI/kt81gKvqPE1LrlQUuS69VoZv4eD5JJZrZDN6HB2a8YUMJOxdLEEDj/fA98j7ad7vk
3yTXVnrUfz3Cia6IRVcIbq1elsemCnpCVlTNYjx+MmUSPAczZ1GWVrFcJG/iWpZfInxmYc0ZJ6CK
LkRUsP9wjAEW1cA4m9sh0lQyKHvOAiQuD3+LtPX7s3JI/sh63GLrqWDY1rwGCVrro82Biq6S8aIU
gv7OBpv2noDTUhr7HttTPHPIXYhjExi1eFtOgumk2lkRwzRN2yVcJg6PxAv/ZrssUxXMDHVgEahL
NqZWI9IYHQyuJqPT+CUeHVVh3kBzKtstGjTlbG0maDawKg1hGTyCrO9nHZxybgRDK2oKhHhUoaIa
/KNbLAAZgO/HeF1KeIh8uKFKJhbARF7mFfdpWZ0kVuIwNR8am0FdRXvPy1rRcCpolaunP4YWdhg2
fzr5aevSMxO15WzmHA36GUtffY4SVjAkamOskMIFo5UYB3gMn7vD2jnGDA2C6pZgrPkTbvWz3UXo
nGs11obuUSaXUOC4Vgt3Ikn4LtCzrQTHEAnukU7RDDmmm1cLhjvG5p4yaIjgsE8iQ+1kkPLpouB/
F4TpGB5dhZiDM+tobYx46dYzyJEDnpCW/NW9ztx50IMQOaOosCjQInnT50Unj7LsrJG+RMPV2KVw
HkXUe6H5N6HRTT+lYgfqsGAQRMFcgtWfma2MP9Nl+VhpACON3oTyolljjDSgbBonqat97CeBQldz
lyn8s9maFDjmFb13/MEp7XL5R6uo7tWjP3ljs4f4dbh6zHYU6dGgsdKqobwr8iEA5LWuk1GDw5eS
3MoNjQxq+dbEosGpNMQNwg1LPo+qMtWDlC8lcn0DFtWZu5W1qYXNdf5F7Po5Gt0TQEp05/O6wp4Q
Czzc1CLCvbqsZaMsz/SwqFgvybh29ZMZ3+rwn3ju0dOWY6QGlLKZpMdri6/fLVVqzVbC5HrBqD/F
gYWV1Hr3qaFMQ0kwzHFI4Mc+cR8Z+Mw0aGgpWtvsRgyOJOTrHItSpfw/4wSBf8GoL5IzQtzooeSi
E/LpIafLYp7kocQADS5jYGyXxrPPNqwOZzHi+8aWhnCmSdLWT29EMwGCoc+Ato8PD2TJRYrkQ6OY
mNulD0lpNBNtC746jCbhUzD7eDkt9f877Jnw/zsw2IX6/RCmR9L3NTDIVBuKMOPyO1epwOef2gny
dbFEki6Y3RG63NGE66twg0nXJAWh3KH6/OifjHlE3wpXPUwLlWXenpzDJuDcApvXcSHfHFN06SK4
f8LWKaDkaCDd3E5n56BbARnntAWa3N/xOTgAZ3W5FCMU3JH8a1CIoHMPqhhpB4IVPYPSkiybvLrr
NpEz1yV0A0eiJME3qNvUqEktJHbMN3mLp1TLhRElpd68HSSRrnu1T53CYJOLHglSPxuBP5YmGTWv
AKvzFzgI66bDDscbl4LF6SJKjcrJ1uOQnuvI6QiLfxd6ih5a0yKCkpsBT/PYd4DJunxafi363UEW
IqALykX2+FKE1dZUgJMMt1FtJKwWX12bDKgh91Dz5Uy9bwPyK9mxET7mg4cqZ9OK5iiroXxEUMyu
eDc5hWjkMVL6B6eDjwRtRF9P0Ji81O+bagR4LDigr8rvpNGeE4C7+bKuNI0hSa+CbYI1YHr5LrPO
ZTQr56DwsuJ51iG1czPZW7adv2TjVHkvNhaVCmLHVFj8Zlt5ZBskiwzCA6PWF867JqpxcIzBAwhU
9EIpaLDlyVrgtL+GR0498epJyH75ThDdOhMAz67dEoB5SEp427l7O+xLENV3v9lrnQR/OUYT20db
jDnzFAUXaG1F8rleMSFcIY4M3xyDW4gJedafa1ZX0poQa+h0EPnzWL9gzqfjBYHt/ErRyE7OBL5Z
8PWuyGucEFflPo28dYEsyIs9nEsmVx6gpaq0+HjZE6ij2byvXuhQ4B4S/VfyXHaVGE5hfSiff/r6
Zo40hFckSDxz6rvV5pk6TCXUH/Q6V6CvwAuVZ+mup3nKgztixMlonTN7cy1LGxjvUF84pPlrXkNM
dMrzMc13q8WpGTWMfaKco67zAu2dGJMoOXAaSA6gSO0TGNcbZRzIs1ME/XS25A7lm3epZxKQqPLy
BH7mQQR87qompUuRDOX23bZfH65Bu6jKdDsWT3Pm34Yc70elXeAuoqOBK/HA7b5qylRVnQQn6BVm
66RZ6ZQFId/8FqOmE7WCywe3890NWD2NKhlkmf+5xGDuB2P9Qhk3Re4oeW69l7KZR5U2MzryjL0t
J5eRri27wkm6vx+1djcmd8KSuz4WtZLmpVFMAt0VC2VvdYZaizfPHMj1/KOoJldNFfff6STWaI0a
qNT1CKEpozFUvLqD8P8WdGIPR0Ezkd5vZil22qpSXoikni83LiVkkFxGj/JOTCwPAIZV4z5qNMpx
k6PyqVAhnFmFTrNqAhoqV3xJqjXO6vVv8++fV8i7FHvAmMZAYBiBb/9FoBsnCK+J1e0O8C1uP3EV
iE745392Ybkm2nRn6Hh0ZmjMsNn8Dwf0cpi/SPHi8GKYKu/TeHfmZKbLZnDUp266yLzOEHOt1yoy
PakJUAPlHSIFHDVYpROGBKqLshutfdSjcrupdxriG0cSJDIvm+2TgPL73rMeyJ6iJT+7BRHc/wk8
J9KkQBQV0TgqEW+s1KQALMhr6qih3uyW4pBciIyiGoAbnFvlNk7Wi9ROfN5L166vs84IgCYMCCwS
93HOm16KILVf5xtTKy/cEDQFdAm4RCPmoYy0wToP8HGl4ZK4F45K00v2ZuQ9aPzswbMj9W4Ahvg2
v00KRH/Ydo67jf21/nDkWUqrC4TxYuAVCu8T1aeQEpzNWrAt1zH0YWOly3f64iLb/AkwPYHgSMpG
yJXp4Jdrfqd4FwNaJl9zl0fAbmQ+x9tJDjbBzD++xzCQp4+YFHAMjt/vh6Na27d0zAHG9L3RIDaR
GKyFTIOEJwgWpdXZj+ZRm7qt7nluJOTbQMMDN/MQz8vl+fsO6je4kHebCeM4Q/Ipwn43sFAh4uvb
jbj2z/jV1hN7/upJ7cV1dHyxHei2501RrcPzKRyGx6t6KcIgBRQuAPvYAV05WAr6SWa77ygywSf2
IGAcGY1EO6LtsKVDB6Ij0lsdmyWGbbKHcf9ZacJyJGP31gVthU1OfcAn4qlRDgmthwk/Oy1fNUU3
8c8PeyGKmcVy5Pbd7phwoLCs5OfgbG7uRbHDec+PvsLEfnVZlA2mVOsHNIslCLNgCVNWlMNjcUgG
CjqZFPxCeqUIG9N0RsW0sAnAvBEgbFsj7X0JXNoGVFkee4VhxhmdwpC0I18ArWYWztVpn6oOLXdK
Tt+S9D/wS3THX8wo7g5jczKSbzK7uCi08e5mGL53YYE3JgFIb8zvnebikTIS9vTt46XPp+d1Jn09
6/O44NYu38OGylRZY2mHHTOUYOYZ1n35CohpJkUpRY9rsNKidWBIF7QGaH3aMym1i4Tke3SniXFH
lRo6KnQ/d7z9oqiVPbwlAS8KWLjiFe+wfwIbOY+/9r63KfGfLAG0Do0gt6savLjQmhltYU9AHiBj
fNt1K+gmAP540QuszibidRIOHOs6qu8P102MRNGlqpQ+3wq6MlejYeShci8aYsCEWCSnBsd/JAdB
sEwrVV6v8+6j8jKT51nki7GrskehMvMuAz2cbPPNZOdVjL+TrydPtV/Tneoa3KaX+aLvbgW9sste
HsddTZnxSU2p1RJm23J4M+XkTzNSYdjsPQ98EnAajOxhK50Sp7FeeQhN0h28ojJ2SPDDAvcAevOd
Y+NPeMd8jHh3vPJJhVgLddC/EdwoRTYCZaW/TSZeG3f+KgwQyGidzgDmHaG4E0UrOnaNYFaqf2ZL
0Or+vHYy2ASe0O0oyPi53ELIpxcj5iXrSzo9pl9NBN5tO+Y1vY+KYqNAMbamFdK8DYTIr6mi9ok6
1537Q8AUTlJpQWqCqgy5FqGJdv++V2yBYLigYX5CzIrscEJlWTHkaJ6yWUM+gGKw29ts9gHeHV9r
FfubQK+KpD9Mfm3HKFwXllQ6VkXbcwSxnubUBtadB3pi37ewKqchyY/MCRQeL+lqsTEDBQS6LLNy
56DyV5cSEX/3v4o3VwwC/ZbUcmXzrhRLiGOwUfaGEY86+IUYLuWl6EOkNGTV+slqbetsmyLbLtIe
/AffJ4JGLp8XW4A7XQBoAV3x63/gd7GPSaqOu0sXup4lIN29OBvhriOmIewJeoGslGEotm0q5Cih
+fJMevIfXjTNVW6fsTBzZkW6w0nKipXnghKOVj5oszGjRe8szBPkT5GQ8pE0+LV+KFg1z++k+6Kc
vHs/3y/zd2YTDA0yFZyn9NZ0uLLBvbjP53fZeBcIwsD37hYvU4X9qv7TVvqpF/xqk6QfMRO7yY/s
Ike1u7BNK0O+mXZN2PKfOIvdRspWSQt+AuPKLD6f9+43I9LD+cWM4Cv91XdN7Mey8YZxXeGHS4d/
w+CdPCIMNKyMI5JyFG+Cbzyt+SlnCBaCYCAkoNYzgOY1bKIgZcWgXZZjnGCjIHKlL9xrOaUPqWRB
TFG0cbI2Sixf3es2yRB8/TOQpOfLjFG1uPyks2rQIL4XxV7fd8lOsmDH1NgF5XSyL8HKUacJjZ1h
6yd8xZ37BAFBV02vp7eZhOxiV0PVxhqLhExjF4LVcfrIB6onkTqd9d8PArnqPn6meSOMPNkPvfr+
i+yBU6iRXlQWrEHCmcgY1SGH64CDrh/6vDZYk818KdocEo1U42W9Gr8g/sok4QPLuh9hqHTdaYyx
41WAH0tu9oN+l68Bux02eCjfeITJkPblqmGXkbEJClt5nL0eRJUjAU11THV+PnD4bm8bIMZJk/rw
fUac8CKO7YSUt4hRqmp90UqunLUf5FLsOaxX6sPDCHxm7MELgm3sJ0rk92uMl6+AmsCR+b5cboqz
muiWUTA+YQKDZFbIcCB7TgEYrsVql5rCg4V/8fYesYTo123MyZZrNxpnTglB8BsPGe+zNUfQzNVe
mENrkAi/9t//kdNewVrNPIoNPHioGNtak1cdBtcpPLOue2P9OFO+pplalJqRqaPROXU+SCTo5e9k
xQmDDQMsvIJy3Ry2RvC/HPJKtZbRWOHI2EDgBtVJ5IZi4c9GkjkVzTCv1zt6MxPLr0c791yAWhqs
lOECag0gQJE+J0E0PFhzN8o43K78pWWj4loErd5kG0p3QYOK/vDqz+NTz1qp2dwrS/rOl35+nYPm
cdhMzQyTpTOSugMVdNGDbSzQ7Mu7jkz0IuPJuAEccZ4SKLdn9FOEFxjRJ5laLZ9BkIAuttdqxphV
Pe+T/9iGAYGw2zuSHksjIt+Kpmkl6pWkhus3qwJQsVria/n1Un8RyEBlNvMlCBuZZKl4D7VpNBJj
P+ICnvnangI0cZ5JS8eyVVqlQ6nkgAP1zMvyRYxE8g44lN8ifwb7ghu5ZaL2RhBi8d6R4iAGtAwp
2V35q3loCg3wB9ksSHUAfu3QOTCzP4vr5qBoyU4I/NEbgzOU96PS1LjuFPj1LHBNz5ICoTwMlNGu
rx5u/QsGQ0G2niDgwEjIxZ5eEoWAJHxReClVAPqb7gVQGtp4CPzhD7rbIgO3KMp6lESD2eJsFxPL
n4AKTmhkb9Ux08eZAuG9UvK9+fRZDdtCzz3DJ9nFGsBQiJuBzQxXKxMeKy3/nxhcVrmMgEcM2ayJ
bwhR9i4VD1UWSG20D6J7y3M4sGbSAHn2cokGLzxXBSE7NhfPhfncPsKqx5EjBHpi9QDGov90Ddbx
RMvL9pNxc9OzcYv8qlz/jRjK+8ehpXur1X+C2A5OZA7ID3qz96U9qwRR/kIPP43QFPzzSbYWONyi
gp9OsI3HZ16WHTg5M28Pv/mklSdDzZ8P4hCvuXBYc5M+BsyA7g9LpX0ptSTCXxGOdSwT48K9l0R3
yFDpZT3jULcVqLR+6Dyv4u7WkU8Q2AcNhDM9YyEHb390Qy72zdDvRJLc4mZLNE0fnEgEwCqhJEJL
KW/sk30hU6Ns8LdDn6Q8AbthLZuMIakVR5PFIsfi7ikczFBfcZYdxfBz84UDFAUWT6Pos2iVIju5
qwM/crsQ2EJB0BC1iMe5B40XyJp5UDcACykch9rqSDvYUccX6OYjsnNNWNBnH6lJNKdi1cBZZZLD
GNJwqDWZP6sScycVO/yiiEQt9AiYTLGIu5reGrtxlkBqAj67stwHO2rnc1HwyTPnVprEhRr8fvQf
keLZHy9kyv9ANOMh/b9t6vAD3FkzcpjHpcwqDwyJy/4dgQjOtp8MBMsrFDhDiNpzuii1DXCv42Ti
XuHjoggkEWqj6vj9uPhbajPqBI7TDVKiNu+6g0paOEU7vsgxyLL4Q6xvkIR7McVHpjBmzMa6HMlU
jS2GqqACBa7wimV8j5goyoq7DuVjXBlXBgHK6YcIkDontAMgVY2MRAVR1VdfTZ1yoS/NCFhiDb9g
a93sad2uR/Ha3WsS1fKQlTbO3yNNhpVAKRv61HVyc86sYor2uyLEDCFP6/32aHuGeH8oxZlu80t3
kayxnXg4x7plCqZhvi1YV7PiK2LZjejMPN1j+zYvO3UkfHnEt05wrccAKiaFr0pUE01206vOVypI
bhqr1QOMz1WVU3ViMJOYlO72qdsQ+zVJi3g0IXNROlrFs4SpwHDL38W0JmHq4S3LkP4vGS44uUOn
QuGtXvzTw1F4/zZ64h/E3wrYVRf/XLVjivg477DY/csPE6LFJIaZHPZT7V//d3Pji2P2+aKjDfp8
TeE6oYcfTGYbFzDL7332HLhwgzSs6uIOeC7I1LXh7kpRPSUFw2STuezQeOGPbiAg68hUXjb6y6ee
b46FHBscUkBQPinLeHNkyITWGOaLt5xdpws1yC5HGbSdnh9v70ki+y0e3BO64hJEkN1tqQ9FvpRz
F1Pn6rw2Ry483iXuZR1/tjr86T2+vk36mgD5ulgE6uLFGp3fEZu/K746q9+fu1rtF5jZSGBzpNvB
6woEQB7TlzDqIZ/ASlsqKl29T46kmyafm/qHFlMHRsfZLs5sgfPIKidCdOZZYFr0AkFmwRdqqcJb
WICuNq0KrwJszze3DfNTOv1gANXQBIzV5RWFL6RPVeerce6NJbmE83VP3F5/GpnVVZXxvTDqEOhJ
mipTHsfEVzhHRL7jipT6EpEzEcDEkAOYA9C7Hv4AvrwwP/I0IL4mpcTwmhsmEXjlizIRRCdOY/zZ
BZVqMu35Y3Fbl1tZ2N7DIT4TMfOLZtTwNPJRKa7TtNiABSCAFEi8uJ5XYbGsG0M32tizu9a5PG3V
z8BWHX/rl1VzJkbcdbFd8BwmSf+X3tnjTywwuNXvqOcTNuiugXILC7UxCRzaq3IIOdi8HC+HRHOd
aHftsXHErih15kWLSWtpfBbTa6F5jxmPsMR7b0GWqD86naYmgAVnOEL0MNmgNkVC/ACgi8ADGubQ
q4IN2VZ05bEf0b1saUVDt3mX21rmK1NqLmAAeudRQRc08th83zdRA0iSbo/Zg7vCEWrxBwURvc8h
s+QUj6HC+Be1x73y07iWdTW8opAsWKY32dfkKweJS3Dd48sXPL57NDyAt7V/ZBJaD52Tym5k0FCm
U7Zt7uDAlepzVYhRqiykc8Q6NDlGrn0o/YpLC8fCQyTx2VSCpCxsEfdAxqkfvSgWBtsZD/cYD/3u
jIp5SA4YfUWitwR7w6vzX5HjAPqruOlxBv+dOhkB3oMTsQxYUWHSlTXhxCWIkcmPMEwNqMEOd5b1
qBf1oPuyQku0Xy94t5u/F+I5fw3y4KCNsCjAWUm87nAEDJdgG4E1YLUdgVBy7b+eioJKSjpUlFm3
PQGh66U9n61a5b8Uv51PZ5Lxwb4OUD8EnbvpHSkP5r/Bw2lNOaCMMDpGziuKTwikddxrbd/NrI4y
Ftg6O/27A39KmY439o9WAP1shIUM9K52I2dsFGbfpiaqXIzcm5S8DXUQYPbghriNwOHPYLlwIpIp
BnXVH2nThfSoJe6es8wlEaDLBr1NkVtxpfSk1MeoVr0mNPqXEiGfL+DjP1moiYOw5cZS5d/VRyxZ
Y5dSSZ8xq7jP7Fl2G03VH4WXBweimcXBFgtHcTIzuo6ma8tnOBsZATZcNb4Y1woBiDFu7iTu8tWA
qSojbqDjOQ4ijti15P35kDGiGoqh19etOJV78j+r4lBmL4M9s4F8G8ZPOdQLyRKMcxKXH3E/0L0L
iSot2dSkTs8lSKobXGQtSeKLr4+I5dZAI3orU6xgHDB2Gzg9fxhyRnSmsuXZ5mch/WtHA6rRHlD/
vKaRSFzRWeVzaEqaNjrm2fdLJ54jvh/7wY9X7xKdr5FFE2m7j9qzNO+bocv2eRT//MC6Mhkv6QUL
VCA8S2XU3BQnnWXx0GVA3d87QMqInKnLFpOu5AJX7iKPl0dNphDlauI98F2GcQaT3yOD+ge9vc6H
WK5iC5RS2yFfAb7Stu/w4fhnI8IOU3mu1ADU0WiE0AgAnRqZAYWlK+14EovakpF8Ou1IiIru9x5z
U+bEfQ3hUN+dXizIlCL0tzA2vcEiEWd2nQv1Oel0tMAzxFUBDEwgQ9RrzgF77pexNS2VN7BgT8lQ
zc0pPQldjR1oKEo/d1/mSEYdai93fenxZteHWYb54/jWagFyD2sH9RAD3yt41NtbgdEc3vEfPQUe
Qq33+Q3AoPekY0BIl6If58op5smAevgm0zaciU+ERMlsB2Q0dlsWuh9zem/N9JgvBk4A3dM3MGVX
OnMzeHTTy0gFjXN1LrIgCqb7kLqqRr+j1lwjoZm0B/K272fHOSNH+Xxnt7PXXQeJHwenPashoui7
6PIX66xxDMyz1OS6SejYQsbReyOkSB49PMRrm0QAUQExCIZtKW/Yz1AhoTaYOGAa7FyC1CXQ8dvS
zjvUz1K3HQ2A0WrcrSDjnx1Uf1WSlQJUHzo02mLxgW0x1LttN7ymQal5hvByXZBIG2qzTs2pYsdS
Sy1EPIGuoCdm3W4pbppYJ7VP1KzIGcronaHnaJdlPIbeoxPndjxxBkVw81o/wED1o38yBJQFPhfN
eLoUXxbXZPLeLypcksPutK1NwRgYeiFLPORsaTDkQPNFZIv9uCcLuoBI5siVgdWjjkfYh82oaF9b
xxQ6Shc8BmFUh3lTIMpEXJbEYd3Ifd4s1IdsfOsjEifEIRYZG3LhMaZYRh+On/rlwONtMSbqjhga
TBnO/8D/HuMmWNMQAvJyA8BgN2dqcRIfi3/EP7pYQzE03J4jCj1ouRItklXgRzTUecy3lhRo1nmN
R3iZnCEknrg77FJ9t0LWs0+9cZADFK4YubsXjz26xbWQXjM12gs9TqSF11eEXYdQEGJS0vsjE3t/
Z7AOOY8f1r5tPVwmQr2OR3NMENLgCrjckv/OY7wB6/bYTm6NkQP2IP3ozp+AvwnDiiFWw/IaCALe
k7+uIHURM0aXXydZEoZlaEeCl31dTXuS69TDszW/BHueyZRu0idxjhSnSt8JGXf1YJ01ZVkfnHH8
rM++RJ6bkd5MwGczdISXZ/MnWotP7NuP0tXSzP0Q0ykCfucuhz/ec7WP4bNeEwTj225Rb/M3A6xi
T7P8BmqbmiwtwXwaRcykd7VK8waY6GidMwJVEWNRTlwjY1fPcqL8pIPZ5VT4uiFHrfJDtaM4W58O
11ilO24tL4RqR2V9nwl6XaIWYa56yhc1EOJ3BFguxVc5726ChrYfnnV/Eae63S29V5nYJ9LzfXkp
+GkWqYxCpYJJeMNIlvI9UxJXV58ksFrXJ8HYEwXiM/BWcW7JoxYvWTu6Yp4ZndiX2+0eArGZ8a5M
jX8F7mgRrb7hY8rwZANXUd8SlHgvB+uw5q3Jopm0SPgKlvO6voR6YIXToGqdxyeCQmJAsmrTmQpj
YGgPTFoSnAJ1iXhC01Eg8xrjcX8+kepZa69p7TwXyKrA/lInxGf3z8Yj1GGhxA9REFOo0TLU890V
ezjWfZOJJgEY0ITEi5TVtDjNsU+0nnDdz90Zg2XcZyKnbWqqz3rwPAWWERYgJidClVhm9Sa6StLT
UJxqPsxcIDclDya6GXGkQPD8LyxYKOiOGLeRScX539H7kQ2buI6BjeTfbYGup7fqaskRqRPxPpIe
7vPKV8CIrvBtNLEiENZKgSv+8F7caF19wy4JtgwFhTZMkVRH8272QyMNCZN5+ohv28Er66T+HR55
fOj7SQ9wixu4CArNwyi6sIM2Js1Ch8c51ldZyJ648KdhXKQyWplzPlNo8advaoGQyol/atCIfkSU
Yq8sNfYVN0QYTqoQKg3qy16FkmwpGfm2ogrliP9AljM3pyK0TvQV2rKdaD35rdWFTciJVOLMIZCR
sJyBSlnBU6YwMmr3EWO6V/k/1rn8wCCRrZJQwZol4GzniaWDLDaVDEy9omPtGbVw9tXmU3TfILOV
2HnkK1vkqBYfSCAcmZ49e9gAl+LQQP+mMtlONobi6op0qjjM1y4y7SaMZYoTe99FS1e0YUY1UKSO
hyMI8/l8zAunDdFIJcv7e137NohudRG9qqmqJ58nr5hjTiA8Dk6hg83vpzm9xjPxO1uqgWz9LgT2
gMxpHM8bPkmfP29/vyyVSi5ql99kafe6Rwe3rNIKShXtzy79fObwAYAJGL4HrokDfV+hMHMRiKeg
ikc6Z4NYJZKM7O+JitC2dmGpnDDPYL3oJGBttnhpKFy+6Rd01lK+R8DuOVFbhUmojRmLIixR+Kkj
ipXfSi6+kjcrdIEaX8khzjBUJJCfQEmf7EosfEyvKoHK1vk/Hvu1WYa8+BTTAoqdIsVEsewOEAHZ
qwqT0VXMfliMJYN4aUzMMYbb5yvzhomabZ/sRbnmXNSN6Ao2O6wERf4fRU1LXzQYCiGBvoKTVymR
q/URdIq1nXKmqqLHIjxFPqu7ZZaQ/nDCdOAzCXaD8SDksS49civ7sOxR7RUBI9/B7f3jOQk1dAAW
bcju6REql2r7Mq9mcZsU1e4711QWf/Iax9iPkBguqulBz2YLWqWrd+3JohCsrfXG/uMrdWWrHro7
c/UFP5B5LAXJNGjYq6WR1eZr/CzfhfHr+du/IjAo6xx3Y8YnZBOR/p9ZzrLXK6ghQLy4kb9V0df8
VqKl6C4AHKU3ZxfNju4rNBK/NkzT7YFq0PRx1rOTFem6cCxBmSKDK+OUfOd0UbzfN694eJjVpQ1u
e1urRkS/iAGVUbZVQqFX2MQ/7tVr1/W12ta/u0LC1xZfAWQ8emTWFCct7k7cUbMg0MUsum9J6lCx
Zui4PvtffBdJtHcCOiZ7/8Q1Iwhd9PI6Wiczc80hIiVAt6liRQ6D3E7QroJOOPIyRyYGwYg++uue
3U2wGYFlhnWUI9k0vb2Xo68VSpuzzn15Et+TOJQDAnkspG/CVU/rDzpklTnXvLwxex5J4LbwJeid
Amq8fIIsBVU77OiJxVGg8OOuBpROlPRi5EmegBicc2Wvnq2ra8lx1dAByQDTchHm/ejpWfOPrJsB
vdTYgWjO0U4MmYBHiilJDyT2tT6+zbY9E8PV/PkK/nlhznLP9s0CJNpcYVQTYrWarImjuZs+eSJd
uHnl7I5GmvLhwO0T0FYYPtrU6TcJjYhoFb8jycr14HNKj62IsTYm7OMU2WinUZDXkvWhT3ALu4/w
5pfRi03wdlJJEa2DiUqmWgsL5gEfq4U/oJOuvZxk3hEGDWfBE/s3IOZBJDPhN1jrySpkVMAgVtRm
KQUTj+9+p935ZSLzBKXmsxVa1L9wNO2rmmlojb3Fs+/E45QnA0nkIEvExmrVpTk1nVv8k2WvTelP
CBQFoaa/o1XXKKUzGtxFCD+ubYods9xZFOgXRPJqC7GVbnA6D5gaqGv78NTzcNbs4jLHSz56bvsA
9Vk9BahHGUe6Av57GJ9atHvFf9VuK6fqprxwtJJdd/cr8bsxQkdJggcyAOz5pU5mb/VlhKMX4Nle
QsAK8d1O59jaix20P30+w3nuuwpXmpb90SJuEzgZC6fe1JI9OgRdhaJKuaFmDwgSDUxcOoGWhRdW
rqLbwmVYDpL81eK4JPZfBmzCYqxmncHWJRZBbSlBAmZ17jeH46UXwPFnzO/WDn8+Ete3XScoiOpS
Fv41O869lrU1pXVOU2hTEvsnqYujdH/ygHXq0kshx80HNwSKowT5D4XIUglKCvHnJgs1QvGVJ2ta
jt3ADmtpnh944phNqVdjurnq9QQ/XfGeyoq57+RdaPK3lJ+i8XpmZhYSi6L9zqUGvk+4EA6H7h7x
OJTQaD7VxG0NbHK7y2c1NBies6U+phT2XCCBIUN6pwMf4I2WeQrl1JhOh91OcfqSkT5vRoNCcJ+S
n7eatFWCmyiDVm+Z0Ss+i7CUe8CMXxYWQXusGpo4nUVkcsTbDu5ggCWrJeemk9OesZmSxM9pU//N
WkxxYCFVS81MgdFEqze5Tg4DXZUf7khntwzhVnZZGRyCcVPQr6p+wnpWKYn7p0p89KRBo2yEOQkB
bJ69eK3DWRLoUPcOSbgWIYoUBR3gI9mWKfkouabIJuvomkWZdlfye//GZuIgohaHNzOUNkUKTxMS
+HPVaZnjRg5aYT120/lzQwqa1ERph1Ve9yMGiHVWeumL0IklBJNyoNaYhI+OqFw95bwHNEfVGTY5
L62scys+CL0NKDH6+1h8+z0ZUluWGsxgC6QGY0tZZ0lF34tqKTveFo+NlsfPooHWJ8Vc4NPq/Nz1
lR3BhcSeqdBR2lYwfQrH6JmmRngynZpYf7qEfKgyC1PDTtMQeP/nKdWLKKT5+LJj7OhvJYEHBvbC
CLRHxbdUVSQcze/PDZX93Vu26w5oa4+vcUMQqPla9xzIjkCX2f7TmCY2twOl1wb1oR4YwlZiSZqe
hq8m2MoObVOBxllu3C4vuCQXjfetm3fXpTYSObp28wkdJCZWlL/sN4kClhCdnuuRqnabOZ4BM1Y3
lDsiCFsxJ1OFF3QA37v05Ct98PQ+OMsNk8yGB9JHRID6KHA1TduVNk8ePGjDJKbmZLUuYMajGA3u
ZxwjMY7ba0MP732QSDoEJyBwftblBfQ+8prEWh/3r+Iw4dLvChPXOdKhmyv2Ur7pCEnrchqc1IPJ
TxflP29Eb9/xt1uE7NHBDz5Tonti8ftbgxRkThgvQgaYS9EwCG05u5eNxfwrmZChTdz0nAO5VvF/
6AbsLkDI0Ot32+n1CnqU5llqcSPNUqLQNwEGbBaZ5UxowGbleXxkzzFO2CGjqJukrxsfVJn9epqq
v677JTP0EQblVs+gflWe/EP4q41pub6AVC09Y3eJvWlnO5WK6BmstV6Efk5pefiAR7Q6j2b/z6pG
BUK45+JMVGBFCmU7JSPNMRBYiC8aGXDkSQVtA/nV/+gspl+WyfeA27muDfPnrPHtOBgABGmKfOAv
gphVwza1j39bcV1LrDXPm0KKCsT/LO1M13PUufxG/NQl030ALKI618MD7hUP0Yli/+vVhYPHgmjG
u59kGvCwKgfSv+XaHvN9J11E4rjPHxsvbA+iymsbSePWNWPAMoTrSKDHcpKptyTYH6DDfK8stE+u
6MZqBc/KrkBMIKLBcErY/qBZ8+WnwcKqGDxQZr+nT4LQSjrxb7HSP7/jJ3J0e3Tx5wLzzaP9YqTS
x85MDCFNGUkI86syUiTnVIBgR2IOLzbkmzIdCJ51DntCjBbHvNSHW0Jugn0/hynB+DE7gWcwcGtD
l295esaaw8I/64hcliFm1Xxj93Aossp56Ih6QtvMmLF2rO69DF1GlTLd1QizWMcOZDZVLu5Eibx1
OmU9RqEtX54SYmDK+eIK6czEZpjmi1NEFitUaUkcdMmJCLvH8WT3ik31XMiGdspIs88+hYf7U06V
t2n1qEGEpMBcDcJrcwLc57TZ1swa9nVYlXOkGr2xsvuYh61stx9pW3fj3NteVB0D8HIwDpoJFkEY
BnDFZ0O+BFj6md8piE58r8iZ4Jw4v2zHPm8MpFRK4IQrBI4HIlW8h15X1jgH9+KQUM50Z7i360uu
QDOu8nNAFr1i4pIobTclXxbxSag4VMjuuzgDurzhBZjmJihnWsYQ8Pxv0s/33Kn2eBpnJDKZq1bM
u3rzA7udukwnsBaL8Yn8J/UVKgNUVkMlDB6FvD7rvBTGAOpSi+uL7H083gzwaqwXkMUtv+bhp0EG
t5uNj7j3+qHj66P8HE8rYtGVW7+o1tIkcybQ8s/oll1v2Aae8PYvVFEfNWNuDI2WJErAuoQ24Vzd
ZEgp9WQXSKNCAtgqMpfw0FHzsyI9sZ/U+AmE4btcRdXB+BxdVhL0B6fEDXyvri2NsTKRRRu2mMMw
U3kmKZjLokfyoTkYHqU8OOo/LM8n7vfW6W/2ZE/F4gRTFuMVt2gmy4mHjvFTImYF2unexCF0t7ZD
qGeTvORXJDnoDpFIjihOSXYBjP0Hxu5EYvbfIO/ObyoqLtENUSrBBnIL6etMb28s19TAhapspIQT
siVAEQlbZLrmR4yXbSS3vNMEhbQDmGLo0EHiH8fpVSilbnPFJWJUW+3oNOj8wU1Zjfa8TllBln/z
g6zWyQOKkqyU6VkCYjrkd1z26s2StsE+zIl5KarVKnX3SCSQHFOIxrPG+PWSpGg12W2jQ0LvhclB
u9aFvMk425kvRJ22No6eUZ9/VtOvn5FPqs90OYfbo90w1VlB5fdXPvJ/v77F4qz3uOfM+5kr9MSz
tLXtWJqN9+8Wem+uIuQZ8RvImANi193aCj1FYj30VQD2XVi8cHrWkiDOgt1xTLXdy78IxyYlx2p7
XSPOLd0o3ER5EFXgwAlaNTfpyondT4ko74TJqdVQWLzFZYizVW1B2tCBxteVSv2+83410rKPXmP2
IMX2O76waj/Ib0Iaq73QU+yaR1XXjVM1jvV5VEsFAy2g3uDFH1aMDoN9H+/crnq0ytk2Gpyff6nG
7L/TUTiV++TCyiQeHj8J7i/a7FjWZ/q3YNfFJ7OdmsIywH1PdnVuBuIwmWMwrLCjmom9Buna+yUw
noPX73si0OIx1PpMDWZI/lXBKsMN00kLj/B/a1zj2hOiPb0qqLH1ywCFQyJjnn7oNlbiwv/8rs/P
Ed1DIugj3EcsUVAIYIklDOAIBHwWh9riwvjOKCCIQPubG8mpHxmk7BmtazD9yroCr+FLxAIOs522
hpgyXdldJLojLtMjSlB9kEhS69rb4a3zhVQQrP5kyxHEhMrr+Jxm/CFzC7hTdw7o3hNxBLmMNfqa
pBOx5mko8V3V9cJrRM55cur3YK3wUcRvb9hn7xBtkgkYD5qqBrJwZlbMpydN9OjqJJOfzAXwDhhV
pMBMAzgc6GHj7CYUrqNAK+vndYL5I3HoBse6ZGyzQlH+V4oQECCroT/txBqJ/QRideJUGEOZAfWQ
RcNHgFDF2RpjCgqlzddMBcsxdwP6SO/5mWQAxsnskH3lCICqfg1TrDOQwu/O0Hz6fuvVc+afY8wG
a1C6O3NPfGk9sAcjkpSATxmOsIFjWsTy6NKOrIHx5LRiSjqNG9pTU0MRBUp+QOELb0Vi4bujLl6M
AbbECiAQmNdBrZoCE4wDeZt6I8vUCfAHqyI60O46tD6hbfztguI36iGDN5uXpSm+RQep3DGpY/kK
JIAlArM5i3ulJB8ftI894WLidYaZGLhKMYZpZHbPRClx7xE/9Xo1JDWDbWar+uq2p6LwbdvP76i0
Rzkil9BWp9Haa8PXDUOH1dVaa1kLzQb0bLEiNdXm8l5Gbm6D25bBR5tufsthWR4ELOWNqdpMayxg
5YWX3iB5bS5GWbhE+Ki4ACYli7Zs8osb9M1/tSBRmMNtf/mjNd5V1tI13tFbeKJy2s5EPHmKtsu3
ZF2FeBn4cNQyUH9tsU+lwVg0fqXN+U3Mx8EEG+NBRy+T69ie740Xx8rmHdPvJhsJInsu/MzH7vST
ywMIf6wFaSPVxVQRDnPjAStGUvwLUtEZxQzEjsNPNoYSYsBobZvagBnbFIxx8bgSxmXeCcnDwvnv
fwML9j8asXkc0WTyWdLDVHNzE6gI7dHtMWCQziIneUKZd868S+Z9eDofHvjbL+VZCVE8VRBGshSl
wR68omiseUnS7JmX4XoN6Y+PrlcpFm3Mt8IoIBQiUuSVnKCY7UEcTBPKdn2s3OT7LWEEh3CQKh3U
CqCbAsvUNzqKVBY1v2VvsV5pC/HVBpc8+SB9mg/rbd8gXldpM26Vm4I7pxZ0/aY7tnnBOVDliDf9
jxkNSGd2jdjyVi0qr3UCThX9tdtPXjNkMRR4tJVrRLAUo0VcmV6Dpkc4zJ3eKTEYhQHJLHyNZIVU
FcIEktuhqTasdHZB3rwfLgJFmYV1DfWFbrjyz4/86KwdeG1OIb6ARmwJLtveMzkgoqKwE7jJg7Nw
WLcDDri7bst09hvzPQvnMtTTDl4KyhAXMefIZDV1w4tms0Ev6uvl3Gvq2PvioYFObp5jKglDRA1F
IOCrF0lTB3SisVJg1T6iYvBzUCqPvghRJAIJmxzogBsyQOy+h9T68CglZQawZd88J+N2OiFyvlOo
AWXprg3GxQsS8P/Y3wat/+77MCJZBz/qeVNamRK8nhnczISRlhY3/UPXNVvG7GhcohGfpLo6I6mg
NX3JD4X6zoEUfRlyVTH+hg2U3t9J+g35toWFOUdAr+CLnXeBBaNAaRxO6SOmJ9PBeML46cHxhqhP
FbaExp6L7InCGTSQC6pv7zukkpkJ1X/ppNVzESYLt0cjY/YOApnzDtgQ7VdjWVE9LYE94BDtA5bd
WKbABW4EAf0sctTQm13AwWW5BKOvi2fRlAVaeS/PjufeKQOIzkK1w7GGf03f3RKcR8YCKPOCB99G
AGdptgc5n0HYa/VAgJ0FaBN2fO7qaY74Hx1KmyAxLuaF9ZKoXoghXMRLO8fwQBq9mnAIDQhDQkIW
WE93R4yZfhISgHRso5HxQmnl1YB93X6kHu216kAK6wVCsdRjJqhbDH76Rw95uRKWnID0xTuFxFxa
ql7JNogcoLNQVhu4Tqmis1bvGIbaau9dZd7P3CI5Fl7rNacbGCNtCyLv/pThINzr2MlnDv3zzliJ
756rPU2UI2pCZddPXNjc8wHt4gNqOHqn2G9wQUJ7eaVnSzDDUhmnF6oN2rVC1NrTRnDIv3/xDjGa
xLamAP1Cuu5CMDBaLpZZVYvRDhQaI7EEnaiXkCDaWZL4b/ENlfgwbGVJsJVGVETg4ypBal/2oxAI
ZT9KygRrhqYJAj7D92mjEuWdDrOH6Cw5BcTBUzMAXNqm5X73BXduf9G3DsjcgOua+3UI6Gso7GeC
dykyRck91fFb0juqehQJq0mDoXqwVavb0l+gp/k7FB7iD5SAkBUUKeSmQuMIyONfUmFgKY0U55Rn
xm8n4vV6dGS7ow9vRT3CjCbk4ZbNLDLZzDXc6RCchnWmECnezmg8ZsnFeqLPbY2KfaSbNyQuY9g8
4hL8e/rbpZhadp8L/O0HwaE6KW/T2jHxxAFb/hQf0oDdGP+/EPj2jtUYhSOz+C1i77BO8WlwaypQ
lS5N05nKOcYEdK5/X89JsTbJH6CvsHNzmrVu0A3sWhbrLPDH1g/wvwlNhjQa92P0qPkrQfHbPQaX
z9/YwPMl8e3qlgjLCa/fiRoRKIivBjpnpBBacokWilhpqJuM/FA0iAGoHd99ZhHvknaW/Hs/jmLn
jGigFWRlIORrqtpj/fPMkMi0eougfrptDgVxlDcw+0Dmyt9a+m1OiVpKc8vORUHNiSP115ft4Avs
QDb/789hRvGciIjbah/+QF5XiIlcjAxQ4relkhslMnrHT7OgyvzIdiVnDnpeR1PrU4DInoSyBzVS
ZTiH7ODFY8IOXPRJQpeVonld3Dvq7o1dbH6ETeEk0l94AbMJgNVRSuf20e12eYxnIB2x86lZwJy/
qESoO4nbERb0QhGlvsLaOGDFSMwMLn5CdhGWd2IadHDgDRg2hTryZm0bq8CSVZ2/oGYzcWvtOGkM
hoij+ta9BzBmOwesvElACNt736bpbZHUFNadka4uO3ymuau7E+xX8uomvL5I3iEwh0nmTYydOMkL
/gqHKGkfXerI4T5vsM3IUC9M0X8c43ArboKw/dbZuo0/RxiH0v8fZk+l5s/RkXaoNT3ariAKITn8
fv5l6ykidpmRjn/lVWFDebS9pbUclqDR4u8yNJyiTmZUum136/Eb0zoLRVzw5squui7eu92zjn/N
qOeV8b2gJUZPQgJqEhLDrIKJPdT8++XmBuyrmH0y8hir4YE7kB//6uBkeRnFlLJ+SnsgXabqkzuQ
R1QQhf691JCABxIHuPwJeGXB8nrYCkkxLTMJCyVAcHROHSbft9h8kHV4An29OXo5tVp/5ELE0o0x
TrkVYHdE792EDvBg0XqItItK5WQKWVB+HjCYMFCVtVP4cKfBUCRRyYZ2uR0+X4JSKJ75kq0egPLQ
FG/6lP98DJOmEx9rnsVPurQFrCOaqpmnckQaBtajItM7d6NhkeEKxHptqV6QIj62q+Km7XJ1cZNh
mE6FmnmuvYf2uBlfYtKvD2uhdiV/ukkkyBqv/S0wcaSm95MRY9EnFPgEa7O2N+P/zjvZA4trvJJy
EMyyRgj9jOqxQ2g2O0W8k/2Rb7NdpJKHTHfLfS1gjmqSR7RI+M1jMcBeFw639qF3Hkv6m5u6hbD3
fj0jynbmlMZ8znAm40mTbHCQZ6s236GcuRKx3rATHFUTO/hNJbTkoRZOcL0dfynOjvuVGNmuOubr
G4FGswUiJQ4sDaP9rHWrK2KUrQBjcwxhzrijSD3q6RS2391+NVG/Ab3M63ftQkJ+DxpMWtp+UsyB
mv+7sczwmTj0v04E+OelUkB/riicvXMR/AXOW0xSumgbcx6Cg7LJh2AErMr8M2M2rzRxlKDKZwsv
AlE5wEsa+ycBaiHWdZ50sbWk72PhS0yLdGnzTmy8OiW0Fsvklcs/OJ0X2BvLTombfV/CslF/OB7Q
31RlefUQrW2BNX3Zp4aoLIBu9np21TR/5hGbAhxhCLkq2FiTdRVJS78wONR1LCATZKe33fYYQ0CD
yRSy1tvn+kcaxs1Yb52ONE3MkqDuO2LvJki96qCJsmdDx4Lc5d7fh0WOOTWhrP/j2NNiwPz65nbf
07XaLt83pS1sAyZhSg6ocA6DSxbnT9rDkJ6pOHgG2n1Tj4/NxogonCZfk0FVhXKlVzbu4zQEueTv
ySqJ91XFFyCl15PYb4MBki1Cexsn4Zn+eQ3vGn2iwjr+unMaoKo+3I9aKOcQ8ZRvF7LnXJB1PObQ
OwC0BXiguXAghJqLsanlm8xXkSUIlk9CjEwrn4vcaZKiQFGQSthgr1Qba9BKMj8OYKLXWvtxlG7V
mC+rHuwEkJu7eDOlGvJ+ls4eLwHTPcSgY4Hz+GX//BQS+RDNbgASotEdShsznk4QZclllnNMuGLL
U+RMPh5FKjk4hayqt5qY+RRVbKpTo9wwviI1q36bW4412g3XpaCbfJybKW3+hj2qBUaaJVxm87Ld
uENvoarKfmhlIhBiw8iWKrT/2gVPVGMfr8JFpLP7xhq9pfsJ06cJzk4/sXRgUHuUaMv1zBxqQMuk
ward7NZRWF4DpFi5vCDQKTyjoW3sPG5eBHrdwG6tpiYdbGUcH/Ai8lCpABpKQEzFwYzJwlasb9/J
JP9DzJ61BcnHBUcnGo40VSaddkOhMimgRyDAKDpS1KHezq7AgEFYrVGZ3wgVbNa3Cfj94Dq1ep96
DPslksvnGITjvgjL4YWGsNPRoPnOHHk2xsD3OShChZycdqBZqHYkI56hIin6orfp2C+fkq4Uww39
57pNttPqfzh6CduILtLgH29kfd/zMnOcEZNSpBkkoEBSQiWkky1J0a5zjCmoTF73j07TchoNDwLN
cHZHYihUiQNVyPK+cAzzJWa30ugRsMcUcsfVFGk7BtpQmIIcFmnBhA3eEBmbgS6hUcf3UqSPQQ9M
u0lrW2UnFuqlyp98ITLqk3rJAVKLpE/9J8AxpsfhhCSbu/KhGVhVteSBXWo5SV/O89pZKl/OyD5g
yfqGtKBn78SI8AS9YENLz6Ouia5PJaJH/ZTUWnDKWKWLitZxckItXncg56/KzKmRkG5kWruiwmuy
mcNZiUi9SCmLbKpNrkNwHG1cZcI69cbBW1WBQNPu48nWRlzVG6CbFbO9ICXwCdYbAAsBRqmiL2L8
jb1FyE673u3Se6avIbMkqXsAi8pinaR+5mpYodaNexj7NUALvNOXbPxfuwrDf83U3jXsBUXc/xue
n3NOoEYs3lMYFHv8bnkNS/bvCAe6nqBgG+Gt0PcSI2MJyXKciOF0JhxrhNOjaJSfNCNDUnVxS5oO
RAAxcs0mXfcZzACdpJxnwTJ2A16RAo/yz8CMrMHbMLODIe5IK/R+ipLCET/Vdj6PqqoWcCq15HUt
KVDNU78WOtxFV2uh4YFGeKKrAtpjMFDEMu7Lfoh6hfgqetyqWSZWIDv9DVw5SboRUBnryytMhAZ+
ecFv+YRLqaof7QayEKQIE4tuPJIameo3m43ZOAw1wC3c1cSz53zAIOzfqPVfA9/T5XJCznIWu07Z
LCsWQIWGw/fDC92eVD5TGE8cwggZEngBgK2P58P4KXkIS4+UpfspYRKrHLffcLHuRTCLxGXL5dkM
BuXMcSf2WdJ8CPPIhCGADIuMonb3Cn1rKJkNyJaAOoLIvZV0qSzMONntSyN4dxghjcOX7qa8b1yw
5x2rdqfYv8tZ01V6Sd7raw+vXV8a7FFPw9zhl2zfe3yQNYgc8QIP71fB63Nwarlw/rgiGQZOAWIw
aWxoQ2Vmk5vTFtqWfUZtDntKFuaxkHDNMkHrPGjSZml5TQYy/z7bfYKvqtX2JDjegap/PjpLCP+i
r9Qoj7Kqs23ypyT1ytbII9g3AC1wZZ0BnEwBcTRzoILqzBacM6jSsJycPHj4uFxFfUFc28K54tJP
uDsCPIDOdB031rBXa1kBgh1pzAlFICPdWfXR8mdEn3LKoycS9FoXWGHjcz6KxJn2oGOUePNHTX1M
aEBH353ugpLweNl5P2FEmcIMsXtlsTcIvPEvl2NuirQ100LTKUnY9dlJ+a6A+1ov6dTBi8ZSecbz
/iREs/Ceykz26g/GBFxYUcB2H26AHbLTh6G+j0tKW8I2ogxXzNArwj6B4OLcS2MY/OJ4hMTRgwfl
gf8Mkz+INuAkP8edDZ5imxVoVkKpymmKm8RVZY6Jl9mcnun5iY5FgSv4UPIpeK8rSLo3obM5O4JF
NHyJD0Hpl6gLjTH3I9Kc8vqezPBN7VhxdSupZ7uWa7FrlbN/T0v5HeVsgd2UEhu9K6X6UQSddfcZ
zuROgMBswsU6ZiSeKrNQbG4n1CvnoJsMYLjXxMj/V6rIISaDCPwPFiUW/8VJ5CUJRoz5oataFDGp
SNlAZw5+yg/aHBgTRR9XxsaDWiGrSWcDLeWMBIKMXrl0dRefYcqIHfKBBYPfI78h7Tx0CqJ69ber
3G7HeC+VLV/vPdZIkNHNmPwxVKL7pwE7BPlXKHOYlv2GLTyky34iCC3tKitBs+fpG0tdH9e7mAs8
uFMTIMdK2laI1U4GXOQls1zSmKry/esCPLApUKgqnw2p8GzBBQ62Y5JAV6BAeT85MQBt42RC48cu
H8kyObb3rYnl2zPEk6O/gGw6ccnfBPQ4KY62DGJmWgpfUgQEEBCgH4zZdZ8CIBzAKzfLfzNWtpCm
CyEfRXG59TX0vwwbF9MR8ZqPZdMq/Lzl4CR3eWxQHzeyfYHztGMKWQCl38/4/ng/npJvtGnBX+aF
iVFMP/utPwmWvtB022Kfa8+hTuBVFVicKylL/YwhJyCXtWVZ2fU0g/hA32sWGOAcxosXPcehRuql
rIMzp+zPf4EnC2pBR28sb7FPTWSQAaLOLViB9Y3g7Yt38KSaCukcSLBN6Hdj2585Ylq+SvSNAPP5
/FnHYHroAS3cKyqRTd9YOlqHPTUH9GNbNffYuVCixCVV+ZkMIs3eHRFo4f91tkzL7rH7m4tINdFV
RCktCHrU0WsKaynXOCwN17AJFY1X9aMSgDE5/Cg0b04FjwwWY6NC9qyUc2W5nHM5qWamDZOTnlt8
5IOLCr9J/Im+DHz6owPHuO9/H1hcO+hzBISMnEFJBxmubk+pGWybzAKipKBrxxzKQj2jpkyZLkvv
Dbli8rTq/8IWWzcehs5mEt8P6RN9UdX909O69r8a+ak1safLcQMAKn4kY64TRGdXQGHaK5Ji6qt4
wEvessapH3N7BuernxI8ZBacP4nbbv1zvfR0axH3RXqWYaqF4iW4BVcBXx9iRs9L8Z616ZzEXJQB
HDsZ+HlWlB8W72JeAb6OPaPGIq95YtaVsewT+sB83AIdhXx68LwKXU3Lu3+3CE1uTu4fkJ2Jp1aY
QTF6Z1DK/XE2VMLIwCoH9eRJcSE6UhSbRWMyKOLD9QaAqyKnXfFJmFy1FngHyWupnjrFlY1d4NQQ
v3OOOjqb75flPJ0kDiPrfHTt/8K3yyfLyeycmbOgqNuRTp0Fqr63n+DTqD8zRewrc05DgXY9DGX6
qsE4I6UzMhVL6pSIfR01//C5ALoyYgZrGB7TxWhoMXm0a6i3SgHifgeyhuWy5g5hKD8hlS7qUySB
0f8JyGfkxjQl6TwC5485Rp3L1Xss4dnFRJRvX0EPJHBh9WiVqFbJnKlH5HWx3/fMpAqlFc2SwD3X
rn4LtvOD5gaPrSUKzeuX0de3bGn1LxRLSRR/r6j2yyVgg1bqZse1YA8LtrIZrgcz52s2zLUIvNSc
YbciXB0C80gXzp9MldnMZLXXdMV0y2IEnE9sBX7r01fr7XB8fdV9TMfpGdzfirGArjae5LrjHFI/
wwcfFiv7YVdEiv1hTQcKJArI2jzsl/M8owzWSRnZ+9NxV4SyGThsKc0IuXePdMcFIHjTpSdi0UX8
Y/QZuWzdRa/WWu6PPsuLdjW7UwCkhkDmp5bncHaBXTYQOB+hsINBqF69IVaH7HUUAIpCwUDKJFcx
poaY4BiKKRPTqvRcZ4neFcYVn62rmFqXVa/F6bgGYzFjb+sfh31FSCHPtG+IVzpg4cnyeGhjg8th
YX2qS7Z+EW7DE/w2nIJAuZ/SDh/f3DlIOrQUQBcPJ2ppG/y1U9xDtwJTHC0ORD78TA6PZRWKpGvE
94PX2NQ1cYDqne++3ZBwCvmtVGdyz15qezDASlIMRqhfSAFSTu23MCyGjIfIISMOsMM6HlZEeAc/
qITvxKc1afwR96qDSaM7LaPPmLx191N0ptDfBCQGXZ8gtoOb8Hp79jvN8Y9EvPMrdRKAw6kgyJsk
emt5eec8dAcA5Htiw1wKulgWl/qnQ/IhDrVVLb05GOBI34POMkVCd8tE0qwAl+tjno6BT0iwc21o
R63iiXdNnKCuunWCcLgHI513Q43M3NRP7pIdou3G851xeBUMhgMlR1uOTs8U6Dear++HScAYFUpf
4rLVDphlg8tnyCADJjIDSE1pqoC5qyo0uJz/t/UU6pIRag4VQz31cmdj/OatYni7e9VDY/KqNf4P
xbe/hfCkaTH5yxoxC6/BHI4yxPTsidHj7ULL5C58oO6XpkV8qHvEWcBuKMt+aJD/LN7JsihlwpGr
KmlXHGVWqNSKC7MW+4ghj0/CdwhHtDH1TVTJ3te+WQFF+5AIiPuV6Dwc+ETIUlSSG6aUOLvHJEkC
ND/GgrSu1s+FvFr9QoGl1ToTyMY6sSkdS1mF+xkkCKtqE70WbTldahoXDrmT2Q8vXC/Vx2fxQfyJ
Pqh5uwXtDEvst6tl0pivdS9FhW2AF1dDQfC2m9aGbW2MM35ebK5oyltCV0WL8iBH42U+wHh2dsam
l0OvdW5Yzyv5iBGhjEm7Zw6gRazzt2FTyRBi6LF7jGiI2hX+600Il8DHo5pZvGwVkPPr7nk7y68f
P0x3ZgcqHnc8de0sY31j+X+tM0DylHOtIYwIFSZZuYrKmsSB670yV6hHL7kchVBB2A8dM5vNsjSw
1EGUeazf4nyUcVMoWXIYou5VfQQfB1Plqv8xv+T6Lr44ydL/rFyfxIVnJgRnbDFo6fopTIp3TiSA
Jn+EXCpWvLVm+HatGQK2pvvwTU4DF1a5hgQE8I5UTa+sNmpBEeoYU1sF8nK/RvAMPJh6eJP3WhdD
d0RXXE+eP54q/sjBGJgS+/4/YMtOUqYvHKxOubmeJLjwZqp+8PqTNPY38pJn+o7nej0o4FyQy+ug
WDuoR35LixZXiXlxumxBG8nGzmRsHl8sVhb4yYXI84IxDv1YCUz2Z0MVObaPZapyz2+rYNf7HKaR
A/lpsin9ZtaRT0LHzEaV6oFubrpN7nJuw64D0YbgJE+5xkzq4ixSqHQ18eXelsxWNv4db1Pql1tl
lELwnOcDr/tnzPIgtlLd9x8cV8Xs4cLYuNaeuSq4j4EdSmEUSy0Q7c1bZYaF8q9iWXKsf3BWXixw
jcTasRNyZBkMKJvrURvl/DWek4gvkTXyGeWM86SPX4xzcAigXU+Qoab/2Qp1H2yfttpuT0sHa90D
fEPcAvqfrP5MTQFpT2Pb6/SCM4PI8Lq9m6Fo50YmDcyXLgX/5+IhcX0xrnh6c2n3K/spa98HFvaW
BlaFwgSmRXTq8fAraGBNbkkIc5S5XF9T22IuEO8PfTLcIyS9HwR5C9Yk2I5pgOtv2bxPgUKaG2ys
RNPJbzE1Qq12qU6PM+tZHAackJVNsZWuRoC7z4J/z2VoSbKeH/x5r0HWMCWUuEXtGz7fYC/ObNzN
Uz8imNMolm5XpHXhgbuOC5Kn2HZuWeuPH6d5XogtLirVEde5CW9X9q589Ny0ekS8ZJ32YiV4WRHc
cc/Zb5pD/CImb38eGXbMJhdPJ1DeHfo3V7kg9M0eZJva8/UckS3ElNb6N6ufVOyxfL/jnMvHVDQB
ym23OdR/HRjZvyYY/9BxqZjtePo7ZVYdwYdZWPrYEbBZtDHM0dHmyr1RmqrXP+4inS8ok7UVBgXj
/mn1e+IEQfYPlgkcZGktNCIqr/akZB2GpVI8aIadg/Yrj/nyCry6KMznYkqgbRQRs2isTjozw70g
mHTVCmdkPWWiHrjUoIoSWBKsrrcjq2LebetH9ZRaMRR56PMK4Uw/6YjCLhP1PasW5WfZwmkERm/L
y6Y=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity WatchEventsCore is
port(
  Data :  in std_logic_vector(71 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(71 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end WatchEventsCore;
architecture beh of WatchEventsCore is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo_sc.WatchEventsCore\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  RdEn: in std_logic;
  WrEn: in std_logic;
  Data : in std_logic_vector(71 downto 0);
  Full: out std_logic;
  Empty: out std_logic;
  Q : out std_logic_vector(71 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_inst: \~fifo_sc.WatchEventsCore\
port map(
  Clk => Clk,
  Reset => Reset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  RdEn => RdEn,
  WrEn => WrEn,
  Data(71 downto 0) => Data(71 downto 0),
  Full => NN_0,
  Empty => NN,
  Q(71 downto 0) => Q(71 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
