--
--Written by GowinSynthesis
--Tool Version "V1.9.9.02"
--Sun Jun  9 23:32:41 2024

--Source file index table:
--file0 "\C:/Users/Dominic/Documents/GitHub/BeebFpga_Dom/src/gowin/gowin_tang_primer25k/src/fifo_sc_top/temp/FIFO_SC/fifo_sc_define.v"
--file1 "\C:/Users/Dominic/Documents/GitHub/BeebFpga_Dom/src/gowin/gowin_tang_primer25k/src/fifo_sc_top/temp/FIFO_SC/fifo_sc_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC/data/edc_sc.v"
--file3 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC/data/fifo_sc.v"
--file4 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC/data/fifo_sc_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
coY8tLeKH/su9UqEmT2f9lzVFCP0z7DijIr8ycjvFFsjU0jywjjohj349LxEeTLljsk9LYL3wmCQ
yGEfnfZ7pm9wA3t40ZxUgqR0S2lurnQdWaTR+fm8YBUAyIwAm2q4GdF4Mm6QfmSRqUafpzjKuSlM
Rmhtj+HSFSEbuqUU+55AnW1vszyX7YF/8v0D/vKZCBrD0cqmo0uM1tdI3Aok5iqP2CvMzV9y3itp
xfcx8HYWyr46rC21RRfBAF7embtXi2KRwLzuJh+V7MzWoaeTHq0X4ME01W29BM2Bo+HhlzVv3Kux
sHGuflw6kKCsDiQjKiYna6P3GNB5MhOozMh2gg==

`protect encoding=(enctype="base64", line_length=76, bytes=13600)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
oiI1tMPjzphHCYNDKvRHqm3RLgZEluPhnzBODxQov7cgx3SCURkvJN0NK4otAGYByiQW3dDqUaWL
8L8eu9BVzWd9KRKQRc3AAeBFR2cZESO6aKTwnucRYIOGjQaFUHzwaZ86mXN+9zprze01qbb6GzRc
tnHmbSyNUuL1XJqAoDOyr6IKcAu2mbgYKsr8UheKwXzRoTJxF88LfJ3YkxirWgtJm6hVAWpX1T2F
cbZo47GgoMkajrzSywlWpOj/wnWisaF/myvyKga3M6Ox/0FRYgLBL0Zk24OrvsL5my9WlrI0mtxp
u11Fjlw9zcKFo4wyBggwjdXVuGbK/GObEzm3V1hO2zH5QACjuHLgx3kxCs0BqPkEg1G76bLulgfz
ZNr2HsXTSLXgUfrPcRTVjPDJVBYAFUCkAagYFelnLax73af9kI1VTLY0GemZ4J7rDDDpgvdHwszo
e29IT49vABSry+bzz2MzPnxjMpuKXtFUlkKlLEKgvUkk4q44DrWZZk3CB+k5P4BUrIcfpzT6LpOJ
D73GKpfN6mhN53+tpzLcbnaXGXJtklzHeEDIXI6VnMAOXeEwr2AM/gUFb5nTzqwku3A+o3r4+os+
JbN2aRcv5XIOEEQ/bqI5WCPxJHo+9umiz8CAdEnZEewSyqPyMFkNO1+P+nNrN4W7yDPGtUXc5h4R
MjB0sM2KerO3zagGy9wF0CJF5p/mkm3lXKYu/pg+lusaj1/qaPIrbjN5drTz3R5FYQpYmjIi4XLx
VEu7kAQ3GxoiLylVZtEL47gf+bCese4nCscvhTw+qYAQusILk0lemxSLDD9v3VwzjRsMHdMZb908
8BR2WQUhctB9OyWrVHCnx+S1vT1Ua9/AvlStZZcap7ftL665ftcF/AFB4SQGI0eOCWQfnMqhxEy6
19Z9g36SMs5nSWDNYv0BhRt4BeTbm17nXkra2/I3D1QBQerZJyNgiK3YIwIITcoqZT/orxGr7XQs
n+GM8KimWp6BRxjn+qi1qrJp9mfd9vo5tmMqapPgw5e5DZ59aFfB2pOn8ujvpSTwCyD+M1F01PEL
ubQDA110iSy2P5E7s3dD6HXsA23tGPrc5iOPLE4Uzai4iq+HtLHMPWfPOrQzIDyOLzdCuQR6y5uK
1PtJ49VptWXU7yNt70Spo5NxXqGHOXb14OO5TfqnZJW1BLX/tgouIiJpzL6QDstOkRSgX1u3Nhgd
10xzWUkcafmZBhi5sGZV2hlQQT5RTRXjxivVqYgg20LDHCb4dmc48SY4eO/ombKSa4XWsDzoOdyq
TJGdCL4iLP5YL7YGXluir9hVxKWxRlPQHMF2c14riDES7zg6Je0h92DamWO4d3oCezT4V9GH7CeG
Y5p1SY0Hx/DqZQq+hpMMGN5mvBPoFaJfTbLgt9qnkCCti1zPROFd4k5BbzOez1QObGG4y0uwyfL/
xQpYwPCpppWwK93a81Hzk23DNfxgDqqScRNhbBJEn+8tRNikmEj5ZnbBdjktpxcvCi8U7BJnJfop
aUv4fOm0b9IfN1x5n42eHwkCdWVJa6ahgYBtfIXy1aHQErUY7h5kLaZwETAbE99XYpTpbYgZUynC
TC4wTgOEYvxCmbLprU6fbnHyO5Nd+8cyvUL9H2+v2iMiDbmvvt9+/tMVq+gl0Nkn1npHgIyjwhd+
U2/mnnp/lJge/2OfBPJ5uL927+l5mF1FaKJgW0o3krrozlZvuJMLefzqzKvPdeP14DbMnsGYxt6P
mBbiTWRvlX06FRhlAUML4sjv8Ip1Yock4uhcXxp+zf6Bqu703iMaqwazUkHrRToXwq5dAzOMdKBl
aL6YE82r5btofsfCyRoeyB24rButfSBthIT90HD4caa4LVdmoY42S+p2TWoU3ehYJo9bkJkdywcm
Dt6p7jw3hpWDAonFiiPubFgNKZ8RIGNawRn2wgw8Q/gMidzuA3bAfWodij1xf8rFqn6KiTqqSc35
VZy0Xf8/4ZmnNI+eO7NlqdTCWMSMpow4gP7crZLYHquYgdE2ltp0lfYcubbllE7SFsf2Dz0Oy8Eg
z1xPhqOXG17/2FI9ccmT6Kv2KqMtSQDeRyjZj+NLs8AOCH4o5dg+7/g+BIMq4bdUYJqvlxm1EtbX
ett0aRlUtholZSB2x60dZXcWRFOpg+HArbSF5FiBFNynBhIJYaPMjEV979osdL3ewrz7Fzo0+XMl
FXyr8nqp4HE4Mv4/c0EMLVQ/MjWyOw78gou8TJvaAQlO42Y/UmuDuS6QeWfqWvX9DvOjNqPUrjOO
qLZwxXy9glV3OLKkYIa+kE6zmMV746jLROg76iOGeoReNflcliokrfmtamUpgXoApGxMJfDc82X9
GZhQAOdbM4UvKPKFynx4ShPpELwHD6wIFWK4JhK0ZaJYTE6QE/98gFaJj8mzgvXJ4CP90bIemjwS
KOPbjcCDZ2yYP2TESBwz6CUZbvTOojbQnKRwJylhZ/AnX1slJQ2KGcxfU8siUeyxas8qDqEp4YMd
q34Nec1gx0gT7/Mk2v9pkrJ2Od0qAhjDfaqpvjUwe8GLAMmHWvgDA5HK2Gq/rfuIY7JxcZBSHScc
VW9Hqejx0MvpuHokla2lWEIFTckRZ330Ohk4TiQVQ/ykEEoH5qGW0KAOn8a/QuDQkHf34thhuUKc
azydMlO0dCO2R6ZJ53KAerzgG2/3y65hPJT7hMQ7UhjMVZ+BeP/xE7No0G/q8igxwxaX0wbZ+bze
YydfxeG0Ki25RMBJ2og8xvV4rwLwRwCxgCfj+mbKj3cMaTPjQT6CNRUkkIGYQh4F/qkQZ/D9FLH+
KWhml8c2XzdJtYHXs7SDx8lW+b8NyqF4xOnsL2kdMQc48/2eEXehpp7DZUG5WPhIAjqC1ssgi2Kq
ZJ+SWZRVTGpdOoRv7JeZHMkVT/TpOT3FCb9/FHJ5tO+xBSdVHmm7Vpix4acHmmbr0+b+yUMHSrBd
pD8J1JVE6nWCfoa/6qcifo4N6apJQyTb8xj4lBiY3AadxmtJgm7WVsNZJFtj91o3qVWco+3IP7JQ
+eyh28YgJWTN5RkR8y6WxgoFk7c7RWwI4RF/JTm12dclJjSgrqa0h6tUeNtAHKi5fAvhLw8m5F0U
R0ESaLFZbE8WrL7WoGKuvxAZcrmXbZijX+SB3JICTCAk5CUcNggp2oj6tCs1NdolxyGMj8WIl/C3
AUtU7w8iz9PahMeWW/yeqfCUhsn7PbwqtfdHqWxBa9WT8zsoHFgCf+q2q0Nf69LeD2Hg8oiR3/kO
4MSuf4JByjtIRmv+aPnlOtIE+g0aCLb5xSqzGU8FdgH9BzxCXoqb3k+xiUbHp4nmvy9S/0UhCYHb
BzxT3U0t5ip27bMn8h+hpVSIxPuZ/XpyASdTlODL8iwVNs147HZJjpz9LIS5FXjzAeLESvmqdntf
gzuTIn3GibPLE/04PXa+I+7+M08YeOZoAmXa0qrtQnL8s6iReJixfukY/fsIPtCWTHytuaf0uYdV
TVRlcP8py8FJo1W3Y89j+1OVAB/n6jWlkwVZjxDcAL3UQdb899ZTX5X+YrRSCZEPYUHXKVvP+F9Y
3jQm/D+W58OA/03CZPKLIvyyymNYnUaF8WE/gQQF4BXdBY1cXi74r2LYmogKXvKrxgFCuxNbjoxX
cBBGaDwupVqLugQ+MtVUWU0eqd1L1wctzJupRXrWXWcEYL9p1VDle0LmL+myOK3K9yg/Ejhpr6A5
KK/C9felRlNA/kUQ12dBdqObsvSdyRWEvAhpmC0d/ZfKFUmI/XR0XlHT4lsGfRW2BxcL3AjgWUpn
ulaDbbQDkkcj0ArxZmod2ehguOhU/eN59UtlKJ4rrhvud9cSnwgPYwX9bpH4bQVDv2JwxzKo7Kxb
SS8YIYF4BX5jxyXHGr6N6gcNf5AjIpvx0UWGyNa1MD7ONUVCXBtuDYDk5sO9f+PeTcTDYlXJoK2X
K7ZA6qAI9u9xm0x2rPKInVniUeyRJXuL7WtWKovKe6xKLduSGyaXgKWwwRhr+WYOKYxptRRN55v6
3rgXKZx4B+GmJUp2eeYBLJI/FZj80W2DqWLW1FFMDxhMR523RcdjTJIWiDxnWthsTUpBQaznV5Zd
jv+lxkU/q5DSJMv/0qujsdMqiD2Q8O1+zwXwRzA6xqrhFP+rbr1rWSd/ctXAvidNOJo5+CBFm3IW
/GAqdw+HF2dUFULbkD6IgBicLwj8tAdHL4coASyyW8ErFbfNGxVduqebq199vYNwx2EXBWogszST
c80zW9Yua1fohHeZR1hjJCitep/0Mi1WFm+XVvgw+Prgps6PxZaP0ia4pP/SpZTMBySRsY4PfZdW
k8F/o9hxuZWIxHpcwQOyggZUCW5TTz9XGBQlu3p7jAc2qwVnjGNVkPavItrZsTJ3evOxKUKx7DfR
uKJmN8h6ShySSXLZH/2DMG8s8RAQic71dWYrOQNydFJzuCelN5F4vRRTz/nG5Z8IgbK0mqEjwaPN
gPBgIv9oCmDGPFsA8GoyXylojhsZLoRcozNJpFPQ86JKhBpoA7aqvvMoFFWZWg1nkernczZKMhpf
BYJXLog52WLpSf7vMZgQPw1hdyeAvfrHmjVLtGEZzOqBYT1gM/6SAqA5EWCv6Z0GOCqDt9H/dD3l
/hjTh2W2lTh9qZjgQK1a/+j+XrN4AjpbpPls7+cQo92fBv+/LLpQQnnjnWNKruStNd15bGHAxA5I
v1FHP8mw8UOHM/gWMHeqt9NKRPfun7I+smgAM6x7iunk6i5hFwb7VcSleHyZaqDOJ8bl3rMQJIoE
J58yhsMw5zDIpMiBVmeyP1i6glx28jY7qpRPe7XfenYgg9lH5n6Xa4BzJ6KaMQaJNDz4UvWWu1H+
m4kBACLAJ1vVpUzjng4nNVazMhN/BBSuS/38WWOl9b8krgxmLLAGX65lVyMKLN7kDlv9HpcQfnm2
m/0xJUdaW5RtM0HlvSoOWruX4HYWXnZ7mfaO1lySGoPzy6FRCPtWRZp3xksqW2k74M6OHYLy4Say
j7yRFo98YiPFW2uJV5XNlZUctOflz2njFxlJBTmqZyfTkp0DSVsmz7iGpbQK2EdQjYzRUgDBGZ0v
6cyWF0bEzSphVlcb0yMjVy0lNnj3nwyjDtCvvDKzfoa7+eHm91ZFjKhYcI6D8nMhhhqxDNF4wY+q
/bxUzD1wyEp/ELZCzIKixEtiXZ+x9hpJIu1G1kaqZ2HdntHNHpCMRW0q8B66xVOOtMvT4dul6ayT
lNNYxRLh21/2onZphsb4ExuVQ3Bw3R1lnDKlAq0YLT+ucce6orRqTap01mDFZqmamudbjHM0Q1rl
XbJTkxth4h7Wb73wUqdKqXmxGraHmKgVtyfFmS1HaHWf8By3cHx0WXZqSpqFGudtSh5Y6AIVGEIx
sGrKTmJHdIn9Ybm16AVRXSJM9IPuWv3loW4JgLLm7D5my8/gzP24i8ENaGyncBW284wNqZmro1Co
5+mOyN1C8TnYmlcn4yY916x+nHNUEPvsMHed8bnZMbkgD3gnhazeK8s762FPFNsY374G8felUqrA
ax5k3wBxRR6E514bx5R4VM6bJEIsQqPCUiQh0WeQX9jJnhBlpZ8jpMwB3VUsCFCZQY91hXa84DyF
in3Y124UfxGH7Zuq6YTtyC9341WMes9B6pGAX6lAcFoBY/yBdvd9ZLwfQ5SyY2qGUsKPwvVRdR/G
3A4WEqL1VnzsPcrYpVojHvNLX6QhM1TcBDfbsCNPKnaEjBT1CaPYd0OX4CtB4dyDtT1KWSMh3oJg
SJb6K8elx7tjJEjtuCbMLfIr614GmB2FFFcb8niuZHkG+a+w7TcnJf+4L6D8PoTjJWj6C//RZFyH
6QDGLIyj/IiTWFsaCIoAe545ZgwlkrpBmtXy1CAuqy8U1aLjjAOAcBp7JUAv1g9NzKcHpT031lXq
8UsX3JJwirptwygiiogFO9VWYPHIOc2aur0XhKbXc64zg1v5r4fOWcEcs8V1JjisLJvXU5IYwHQL
Ax9sB0i9VWRccmsf8/aD+W85h3PqlB63XzhhtcS9aBaPeADp64TKJgQF/LHI6hWRQYqCnXzDKVzw
GYrS4MlIgeDrAAgrA3fxAxz4veZPqqZbb6GJY88SWvve4kyBzSHMC2If2Fn9IHHSbeVQ54Y9YE3b
1SgiWN1sR/YPSXKBmEBVWc8+R2pLSxSPMYH64sZtVkn0r81A5zx/8s8/vDe9Bll1LawOtCmmYnrl
UG30CcAHY5FZBx5K109D2Hzc7vnhA4kTZiOea185aV7KreujnilsuivwmctZH4/sPCty9m9ESkr2
L8q0iCuYF5ayBJgYZdUasDTNuMp5YWXG5TaPdJ89pvqpo8M0+Pp7D9X3BfJ1WufUYYsuLfP0MXCs
AQHmzTESEIYeYKZLQmkCotH/Q0z1z2/m0K4Nfud5+Jc6n+TYZCHGbWaNY1XGU3a1X3ZOYU/KhF6E
KiPSdh+ZQ7N8u5PbNPitjuX3YpM+gPTg4JUuWv90q5G/I4rW7r1r5j7x3I6CSgJlkFU6nmHJU5r7
zw29vPQhU8bOjMcV8/SQwWkXiUoRWtQTrNki/ORSfEtbekdJeotwYVxcK+XYpVuCNsXRyDmBwGq6
ia4bStPpBvr3K5aqs/ebpuZZi7CMgRfaB/oKedQTPzzBZGzk3p9jouzJHg1v9+UcqtLpIoBDAVKk
x1HldZivynoc5B1WMJ3v4mGaCpCRRozG3Ihp4hGsgFp+MMmU6Pwk7HFx6TxJy0VTDWHikSViYu1x
TndzXs//EyyqwakNnj7j2rXJlRGP+GMCJ372svOg/wf6DSw4nfotUwggS9CgNvY+DlDTVW+QoneL
EkFLBsJ/RNI2v4p/U4bsJRI9siGdQ2VeHfRyCfnvwSRQrW+BLT7g1JZAmIFtu60cW1ev92GVqCO9
uBdlHez+QiE0F9ETKTxQ2D36Ar3qvCFHYgxRNWBKarMY+ydw8ZZVtzZcNAg8S6MKMwFfDpkqtTpN
toe8egOf79PZIL6vkGuqhw7JwjcayFzhpZ+iwpyZ2y6sDJifHQB5kEEnKb6ev+e7nSeQXyPggSyy
WCvSmDZ3mU8QKny2ywe8oJrl8vgDvu66Sm7fHbvCmsThMpH0m0w22l6JTKm5neMO5XtMfy2Os1Mi
vY3YhhPKMw9a9poeFcJ5sHPqjXeVXMsv7OGOyDuO5xiwTbIMg9C9TDP9QESNg0sVmIV1GJTD004i
yUqpTZrTLCWlapvRGuAZE1iQOFJpFunK93q4hIBacyTZN0E1ZZvDRgrwaHzSbotaqdECxA/NZIXL
wbOfN+6rnQ7yl0ICLsREnBctjejqQXGzitFr2S10Fm90sWcMKP9Y9kUfOx5O/5LBfIiB4rof/Jpa
IbM/cOmTMdbYwDM2xvLsLXy6cYMRiJlWpnIo7MW2qSc336W7tDuu66loDbaVeZHiAiKhBSMA5QQt
zO0rEeI8L7oYXxfzlpFQQHsiT/bwiRf0vla15lFbzWpSxBzhpypmquGJJ4wloSsJrOTcD/YJ3Dmr
bZZ6QmOcom+N4Rp/ml8wB+hQOKBCsGaRMA/8lfmW23tngNDop3XXQfUudWFfYm3WScxtQ1APy7cX
x/oJ3DuAX0Nsf76gmqYUCfNGIJyYO/vMfqWYKARgfvHj+r/5B397ojfkGkDxfafzGtxwWUgmru6+
W3i0mO+LRiqStyOTq8eCErfPeZdq3WGl0qxnikESdAtm5IzZ5VQvkmOp9aBlMGE1AsBk5woOvVjC
S2G8j8ZMwEfwAaJp+p8MGQbFxjlQ06GQffgVA3Tkg0ltPdPHseNThu2JIX+T9MklIRIlhYQeqGEb
qib441Tk16PHHstMTGh7zrfZwStaP/6cudYACe04ZwGtSOuVzuQ3QGg7cR1ChxxwNb7J7+tyLmad
PvIAFHKGsSaARmbhhe01BpqA/Bz/psHuewgwMyrhH0hVSJsuvEvVieKuD+fY5AOwP3x9OjSaavKN
PCTj1TIDN4/qgXSC101uMsps4Byhqh4r1mT5gk23Ucsm/mSYOjdB5chQAyCnJ+RDbWT08MCgwvEP
39B49ZAP6/S+O0L/pOv2aOo0YCofRygdfjlRK3f6k15aau6tgViNSo3pEdWUdnxOuABHppFZ5sEG
K5fFXUO7FIoI683Untyl7hNakKt/UZLRRkiZBWxZjrRRrDqAs6lr6pjdxFVGMeloZCYaPE2QDWAw
t4am8RY4LFXEf68N9UK9tc4aBW3Owvk9JOjSMjlml2b6g6RMfN4h7fqEGqzwLj3hnHLFQzy52SNe
xkT3ry2hiYDxdY9ssTKENTh8OXpp1K7eIyE8qD92Oc8Anq5pxWIMLQFmryiupF8YZqECyd7fw+ip
voiSx9IsVUz5Nt3WgGeYPFJSXRJEfYhdFYNi34wZXLAdUEBchxSTGGuCe0eL1Ilnn/ZZEu2AuyLQ
6WgwK9XiWzDURop3BkhAyNfGcATUf9STRsaTD6NyFAl+QTrosNpj0Lldyq+8jG03rICNJUI6humc
3cazOopL+fnbqMnD2RgJS6m94fKM7Qi/xDRZZuxZ6GG6Cu+F2k91xulk+puh/wMeErVjX+pit+yJ
MvvvM5OCaQXKkIdyxIBOUAxRVje0Q7asX3AAKf5VD8ZSLfIaxqvOnJgjjZqR2XgRV0U4oX/8twx7
FNlEop/7bxS85WxIU+yqA6IjxG75w4w0IT/YUGNPohQ/Hhc3+UhzZjoY/XZ7/hkVq1X+1XUvnWay
XfXQBIyYxRRHbmXFI+WaicBdRM/wlwW7ZHYGIuao4jxWJQpfTrx/mC20mrSrm8BR1mYLbQJRVIi9
HS6helSZ36MCffxG00I987ghIwC4UFgJlKAwExBwek/vT/Nssd6OtwlxIR4GEODKfGrAbvczytbL
i3H7aRdV0Cbec6lj1n9u23e8TM//eOIV1k+h4y/Q2MV3/av+pXkNzB+4dwonUuc/7AzSm1Na/XAC
AUvfMhV1o6FckHH62HW49FSuL7fhUVuGrjFe9cCadNDYDbzF3kC0Ezzs74sr5lM2CY7hjj63y1J6
+NDUzsv8vE6ttwew2e4XNxAq5I51h5eQP9aUrNMpZJGlgZ5igfjVJRGxQJevKghr+QcNYOjuGxTr
Q/BKb4BToDrDWxhosydZdSjNec0XIUn4fWawuO5e4vS8mLUqnFsFOmnSSZZexRuBpPecIu0bAQSZ
ew8yiJh9kPr/H36rikdZnmjRJqJWP9Tp67wJxtFt9mgpNy4/wIdN5/H5E1bAzzQ5VzmxGdVi2hO4
XZvHAu/iQKm8nMlW7aR0wmxjjltWcVPYKtTsGkajspwWVxo1tac3LyW4q9yvj48txiE+TF5vd7EE
29xCQGzfC/zA+FFLuIdmAHFgARDPrizSJe+EN2QaS3mLeh3boM276DeA5jiUclIKMKHAz39WTtfY
CS8m7/Md4Yhsechhzkdnu5OvSBGlsVjEWlTFnkv95dYQ+uGyqdbPh4+dgWFsZCUXrk8KM8jk7NPJ
5lv/8jht5ikO08PiNGw+PbVflyB0OFe+285CGxV/9FppjUWP6sdyqK8bY3SAx7dW3f5kLYAHj+vn
647PDF50ZfDfkhznJixApc/619NFrW2mQe7QPinwhLG2NgVCz15mIr+tAqb9w9Jcp50uUgPB+I4k
ftNRkNA1KO8Usxqf85ie6JXGHZvF/rTOVyegYNYS+Hio82MF4WIExgxULNb1cdKIpDFiR9Z7ZaS7
Na7ZOFJTGZcQsKr+KZVJ2vzys4Ocrb/4rUUNC+drfz6d7zdZ+4WUciNPxlRUYg8An1Ugfp6ENA/k
YaetEYmmTULoldq8IhugTpZnQs0iehPJwA+JJ7mKjMFGOrtV+ELCc7rpSJsJEB2jRlW+fw19da5z
pgUI1zsXjz1aMgkPnWbyck2GPV15s+IwqzSUj3vJAE6ULFrsuZ1cFRhKv4AEZkrtS5F98qZEqzKA
Dj8iRXRe9syUtaBkEXB8/0o2Ro0RqQOxOk74QG4hRVqcUKC1xy3nq3B8FTVMlA//0KEEAqib48fg
3cpL8mkkaAKziAJWapTRgYo+DA1cb/Lhnp5jQKYKUqDkpZ554g2vIULeGDaSCK6d/0FhA1zGJEwQ
XwmFOxlSPjOCYO4a/kj+MWIGCDKkt2CuACcJM4JWWHjGjTdp7TVF6xXCO7l2ik1eC/W2GifvCq76
B0R1MpfBQrV1KskpdtF36pzuyQ6VHaHiKOgqtQ13e3fJSSYgOJt429CryPEhlw/vrt/P16ifVQvA
YBH4nP7qj06vcCnaUp6jTtJXpMiLjGdXZiA8aq5+4vAEIDx9YTvW1g+WCMpYpmRB0KjNjd9EYu+e
g/fSZ71zloMPA5v4/s9MSVVPwlI2VMCVK5Tln8B4k021kTC6H97pfqnoIcREzctUO/lhK0ztou8h
BWsEU849EdQfsgTslZdCGweBoG9Z4+trW2+8iJtopat+gMQ3eTIGc7Jv2dOz6TomTacgWtZtAQ/E
UlTJnbFTpUa4so7NxWn4rdaNXuBv7+uLw++Qnb9q6K0QIyY5+NrmtN1/lgCee/P2bPhBhiU+xUnf
7QupjXPiPjRdigMKKGP3kvCpPwx/kcva/eZbDpIV//M2QSFozlIGB9T+AGerht8uUaZb/zmMUeTy
2plAM8x5rHM50heGOHtm+5ApT+mz+TxlUppA704mqJFdbpJbnLCEVNZ+bWmcRx57F5x60DEg02G/
0qWH9wkBcfPbYBPiXargUgZn79eBmVLWMOp1deOIyLBe6msILRfnnxlL/aFMTtIXyLXISPoug6YY
v/FntSI61PGrG1EGv3UT9MuKHVZ220f5IJutFSyxNJuIgCD5qQZ3Gk0hu0xiia0HJGkihFO88MCS
76dJR/iq2GGXJzyJVQ5UvD5V2s/9M8SxT8G/ruULxg3eiJVlfX73UaAYI49Tpwr8Q/4EG7NkMQ/U
2MEbuNxexEvC6n1VTOtpgPHybd1RoogbjQZfY+VnR+LWYMdx+V/1qG5a/t02vV45qpc1RbATsgSA
GgXrothDkg5Pt3xyDysZTh4zOpauVYVIfgaimxbpkrzJgMzoLPwN7Rl+AnR1xmnve61qVMnpou4s
PrF2OrpFvzKrMF/ycuQj38S/oqDMBJXN/hlk8KPikiqyjGvnTyr7AfMUjQy9hkWXybCkWF2Q8mwP
HSKfWcPWX5R0sMh3X3zSCUzYF4rykP3IfJmEVEIJbuPi/b5NjK1aVXM9QGg9Ig1QT3ei53HJWOr0
jIZY30n79H/yTU/oCvp9PkG0PdYeTNYMWbr5ayUQgyNBp7Y4M7FQdl2/7+AvOJ7kOVXfIx6SkvNp
g02jlLf/e2s1qnY0Zx7NiPsGpjDP0iSUX4vBoi5F9S3zqFq9eawx3prxYgon+FuZsPFgL2KeCkGm
BZ388BGUdx/kfZzCXrKUKsD7wDXv3zlR5oSXjHI8kkgyfx36lfwoyD/fjp2iea2e9tmZDFKiw0ca
fHqcB+kf0B7JyRiPau49F+IG8UFPWs71fOOP8QJKwE+43OkKJr4O+H2cskh0sta4GBmfjB4E73R6
xwWPWFnmWAxXtrtRucmg317/dpid+mjkKHDQsa3iTWgWg646fPEinLwwmJIt63Hf3mNOjjE9AcrX
ZXZnasJ/+ek8gfRu6mYq1wOCsSrAq+YnrL1GRf+2ghxn3ggWUk3ATU6gs911WTm9FeuLR/ieiP85
w0KxUiir2mskFj+hUCCOfuIC14QqvmZ5WcF14odNLLPiLwu48LvgQmeRQp12fNQGpxQjMkYZy1it
nkBVuxsmlaDuHFKDdF1TcaU7TNVPCO/tybl1O9Sp4tceD1QSoWVNLsdEvkVHrkCpmq9g3clC+IZS
ZuXUUB3DqxPqAOcWW5zx8xqA/bepoQWZ66fxYSySFNoqbUqlx5aOErzNgiDVrxaV/taDG23MuIYs
hyR01UH7T+jJp4+Yxrei8C2Z+NmblMQErjijklBOO9RT39oJeu0lK0IFPMb0iRIr3HJiZbg5L7Jc
/b3P83XHDfBP0ANMyolyUpGlSZE3PrZ2ojy9yQWJanEGvShsElzgq5Als6+K+UtVZmW2EAsqCGsb
0TGVWuVRs2m04VMaheqIHkws/K2dmm046PLI8BtdvcA3MAZ5gGv03eWdD9E8SyI56jIfRKVKyUAJ
Pv0AIR53JHCgzXXr48/DgHPoFTziC9S6IJnqUp6DxpBhGOueFMqLQKhL/H1Avb45qNeRVEsEAVVp
REUJ71GMTl99IcYjkyK8mw4F4uqfBlrjVNEFUY2WazpcbdOFtdpj8pcIfZjARPp6+ZZOkQsJgmco
XkPfUnD4+BKXVONRdhN05kFQSaUVIB9UY3LGLEK2Jw7raUB4yz2FuzmaWjs3nYLXPGcdwdW+hZYz
qdbWccdtPeBP0SnWfho40kvAA/jeQ/jKjNqogN8zd54N6uXswxJ0FsSM6YoF0nD5l0eSdCHmDkpI
+V+aMiCzprb8Yiw3rdnIV9BhDa1tbTl/xziP4C6e9EcmSj166lBC8v2RgGFyjmrX8/MSJyE5CmmT
W9NBARuSP0bbGs6/C4dF7W8ATdtD19tUrovcPsdWVwxqdq936tvbJFhosXhq3zccfgq+XwffmIqu
ipbH6R4FdwASv62mJfbKQ04BBQCoEDKivAr0S4vNajSHR8SMRgT+aXsXlN7E9foj6AkhBRkSkzE3
oXIK8ikyDfTIcDO1ZBAFzaMb+G1kZ7a/lUGviV4rBNTXtn4eVTqW2q73PndLQMDSPVgWLSmqXpnO
EBVD5H08fEcQjpAuDfPLlGrJMoGH7ug/vzx0QcgFOrpNeeVhDCZBqcP4Itc1vW3wxQAOD7k+gOmk
OBgXf8CN2+b4eROz0e1wjTLbn1ABjwtH30A5g2YMPIqGRqMrCXnvWqT2IiFtxiD5jHKcFRKTpx/A
FH7OCGEdoIDuWZ6UOEYsOAuJ3wZmqx8hKgi2Lk3/rI4AxTdC6d12Ydx61YiqvX9J+KzL1tLHV7M5
WKJ96BwVA/ZW3d4TigsaCwD2BUInzobCnhBueWiK3a2uhPdRNU+qR1f1Tc+VBBsowGAd7czcHY4R
geZscMYyjNUYRAlI/cpugcWTt7rqD19sCY3wAjeBWY1gjy3Bw+UzyJl2dr4oI1LCXlmNcKmLe5v5
tVmypbvmX0K6CqhryNwn6aw5jpyUCZRu3SSTuNG43iyiu3Z6Jv752sM85NMgdtO/tLLCBfJPEMB+
QdwfPPb0ZwBfseuDebw7GWWG4qvmdgmZPDm+VArasF1D9DpuLv/fwlVWiuokfzx5+ZtZi3D0ja/t
qp/LKzSkqxSe++WeCBKGVR0W03chSTB3PyNOYoPKfe1tBSmNcMIuvhHHVl7b7Gdbqu/EzzFie3vK
ibO7HlCiIUJBDEaX4iBmabKYdjhrTslR3HUAak0h5UpqCa6bEbaEw9nNu8bT+mYlrvSn3iGEgeGI
mPHFZUllx1yrbje7YEsN0E1c14jonwLG9QAEQASXfK/4IvMsaJ/OcH+9JH4g0um0W/GINYwjjZK4
g8OZQVMafC0TEqvDriwWL3j3vMoRNSMX/veEou9cCLo9vWvSY6s8m6up5RHyPQdSZtQHjm7dWx5E
FfQtvMNzv02uaY3IycXr2mDFSHr4D9aLSxNhiHIcv3BloPIBO91tObOWm/lZz3Q1aaqrp8lpR2KN
ui4vu/nNO8rc4mLD7lBnhCQCYLNnhJwIQg4j8G6v7UQsJf/46QGl+abFLipYPLERYH0EsvdyetIF
UluYLfkHdVmge50zJjAccbhj5+TaUDm7pr/IHQRfMfrhjipaerz72XAs8R0roXXgh/JDuqzaC8A2
GB3vjUbOG9xCtbDCFKfTvcOusoOYQ26l3AycqdDNydo+tQNBJJpNTI5XFARUmhySvvtpYppcxV8r
D0n7v8BqJxfInDBWTArpz5tALat8n/EzNX1Xh+sXvFx/yK450QYDPZZhRJGYKeW2mNhKBrF/4eq8
w3eaJ/e6Ap4LgsVgROLhuGi8CQsw/1N6MdhJ2xzEJ1t/lHGpplObG+MbtjDbEy1t37DIfAjY05WV
Ec9b0sk1VdQehYp+VDFb00+gvT0ERNDcAy9nmhv5+TApwxvhAx/U7VlT/QUOOTwzqY5KXkBU9BA4
Lp5LgNh/AknNvXMXgZfmbUWAkx5zIp6evBB/AnuT0fbWHo1KjTgWccl3eDO2q6PEzQ1v1tPFu7kz
0PsgvVBkjPW7lrtg5F1812/jobFfCV9TYi0zxDbjY6KWFPJe5l0a9VQCi4R4t59dlhb4s67rFfan
/lEOO3lgzCXfI9mU2hzA/2rU1HnGg1+9P7uUTFaratKkmEf9+WO9WiPM8KOl0kXNzorZHOG2eFa8
xVTwX6wWaL4289apj5Cazs52+CgPF9v+gG7k3jpcVcAvXf14Ge1d/y6fNtQHl36Wql+RO3CRyKYQ
ttOQlkyF9cqAU3ZUzgBDYeIBy37F1CSvwVp/9Ct86t1nBcppq29KFxYSAxKIR9hcvDofVnf2lBzH
ovK0YwoM3ncA9Tia2jLYGHhdHUIa9wd8rRKbJ6rAqc/FyhGNad/WL88bp5zgoY11TpIIHwlTfgZa
uEndcOlq4a3EIV25Uy8Fz3xUhupL7TrOyNhf7gJJAJTKo0mbMDGW6EbRPK/8TUGKUGcspgMBOcGF
8SC572RQxSkDbC2NmBUw2vzkfIUQQvqTqT6HYH1aDVomlqYGoOaYbJ9vNU18Srp0oGoHQgvC0zCK
SIclVV5iKKScIzA20cQoz0lyJe1cmvtITtGVXrkvthvGy2+picHwiRsqABE3ALL2ZVmRm6V8lYq2
JLLBQBgYV/ijtJ+ksSnN2/O01BitFvs3XA7B4uv+7zAfN804un0Ld9otmSXkarN75uoZxKAFl829
Wg3vH+UEdaBIT4CGVw1Z5kcN/f4ucOWXFFSo1hdQIYUD9WcrbhpXoyM7c/nAldB44jjUjDDX/woR
XPsp0Qc6yD5pF6Ahk4rgNQxZvzz9xlVKK+jcTYBGNAWNeZSq6T5RddoEY4Jp61t/uo42Wp2374dA
MRTvnrdYJSnjVQDGFssGkTOoZX1kLJThcLdgDUaF689NxBuTdcnn6qFedttInOhzBTVq1lhrYCq5
HZUYlkjD+3CKCJhK+t+b5MeupA6MEBlGTICNQdUviygkYXePTJM8kPOj8sHPBpmPFMMb6AImEh0U
gcYMJNFTp8c+vZMKirCTd2QK2ZVABjO8BtBMwIVIJorTpFu2eXgOLf/y/iftqQ6hvr/D7kztr0Fl
Hdomj6gbg6FjGHQCtUI7n2k3G5iBsxoF6ZrDlCdTupWDe1AT6nS/VD0DSZILyUyyc4czixcH78FO
iLdp5Cpl8LCE8T1sKcWrkf3JupxIgC+pnSEwP2zdxAOciApIOjqnjGBY3ZA78jBlFTFo5Iqlv2z1
DcBbUF8zBpiBWavl2Cza7VbMnytlhUZ3LPAY3pX0z546I6eF3MqMsOr5wbv6p6DrxD6EDV1AkDdK
ULcZ3lnX6ckszesxTAC/4ExFmfzCo/Ch+1h7FjgQ6vjWy1lo+XGJqj5PoWFINxqEAcoCb+3W1RTG
OEjWflCaam//q7P2rn6t7LVEIwUFt/hxEXDSQjpk7wxdhqjI+Dh9HL5LLrAIO/OeYVfOlNoh5uud
0gw9zXKkIHbPx1c4OddLkAVmVkAiE3Zi9LlIgT+rIDrkq7AhT8PKIIeC4c8XZABNEtOLutF2Pdrw
jGch213+mq4ae4nZTryXzcg4nmxTPQ6nZYV9LTRtuR42Lc9UwslGQ71fDbBhu7axSb7yU3w/6Y7I
ZbXFxqSRCgy6R2L0TwL3oBJf8PiYT/vQ08SzTIi55xSCmjOQ44Qrqekt8zCUsAhFx8OM4MkXOr3n
djCSnF97ROiQzAUuV4bL4SGnzdXwlZN99JIlK0sg/t1wyGrLNdXODABEYNOk/sT5MvJRQk+tvTxU
KXWXEpZMh1nXtNyzNTtXi4ZnSb24AXBfrSk7JEXXr9FHrbmo+2vaEEmVaDoprRl0TGI9SQyhyx9C
6XAAA6SzDex5e5VN60eEtlCYDIKGPkGQOscswFEl2JnU8SFy2VD/AfBdgjoBtJLHq69IPU7BfcAn
ehchxqKg+uwzZKh3xE0NqWk3lTMUjzXnrnkJNUSYd+H1QfH7A5vxuXjJRl0DdfyhnzFGnQuxudDv
0e8dLz6odxkbuGO1I6NY7gxoXqW//G67ibsm1bjiroQxp6kEwHd2FYe9OEXzIJg3NFnOzxwKE/w+
HIyG6D6Aq0rdnXH/T+STSfk+Qyx/uLW18WJCDS0cJKQkPby29MLGkCJ8jb4VonzOurdXIgMjoSEh
Arcc6tWQvbO3rNw9h2qU/7gLvH3FAGhosOhF9MGkFgIHvIx4DeYbNNsOqpnBY9kRuvkEr5g2EDiC
hDBw/MXmo2mIOpgUlC9ccQzGbYXKC7OgTubbnFYKruOXMPyjc1VtzQZmg1PAU6AqPTXU8rftO/GU
ybs2qsamAzFymyqc//CYcr8WcFIYVt88tYClE71nnaDl93rJJauYEbVPB3QoSlPalTByBW/QfnHJ
rRkQzSqFoS5b3Q1UcSb+5CF9ESmzqKPsInL4/jzIF40+89gJq1EwHvjwQa58TTdeNxEzShLtvJJ1
9TEEV//Vkpw+LXBbDCDlLU64G0Zr/YrGXfD4yPZr7QYFx4M+F5iqkSW0f8wZ+rAOW5jQLr1/4vV+
1Tu9cb2vQSA0IfHsSfAgTtHwwphoJSeB+fwsRkjeINfq7POPhsjmU8DC+p+meRZcHjnPuRYZW+wU
WYm2xdkX/cW1lGvbdfjB/C4I9Lv2x+K+QsC6/qThXr28TaZbZ5Poo0lFXRmzY62YHMYRJy0Tc97k
1O4yxR/bNLaJjtELTqxhcgfTS0Vw19dUhzaJMK+59tR1ED+vqFkANwDCZiJEY50l2h5eLVAVm4e1
q6RK/puwDPjBCpszeDu8sOMSaCxAbGFTjsDMJPcju4LkSOtaMD5spN26qvu+n2673ueOfDIoxmxM
cTQPhuV7svcifQTB8vMkXq1a3QVVT2xT6gPI3dfADxXKdtb47+7Apf84UYUgyjotozG1D/K0lgU0
EXLscll0fCR363FOPHf/rU6mViF/LfEUr+tPln23r7loyY0nf5cVFmQxjVTT+0fJxD3adggDK4uc
mR7jji3U6jlCssHOczpYxEdLnxOQlTtU5whqjbfLcn8c6Uo06Fd8FWM1hcMYJ56zdxejiS4h2JC3
VNSj6i+QfKYDiwrAPDSNCoN7ktj43PSpuxtkrFlN0EIrkc+GFzPIBXVGNFej2gKQg+OPGLmIw0H3
Xw//vECe2H3atEuh53EAqtgjNzdlHx5jZl4PiSbV+nkh/fcd8/zFFLnbnwFy1iBLKfFzSIbHLP6Y
eBKTkyjImbNQ9oaO/TFGYyC1DFZQwjxhHGywzE4N/OSbhbqYLfQark5G8uVK8XMkzBRk8wBrjiLT
PTDn2QyBWV6duy00v+a1HBGlBslOLcfhN/FHRCZ9NrnGu7YmlXnjrH7xx2XBe3PeAestVplTcW2w
sjvEa9MnpcDSHTXXbPBm8MS/fLv91u8DsG7Ois60vm16D0zMkZjeciizVKJa10uXV2cVDspkbhuB
uZU4Z74pfyGBiBrL5IQByZRX1ImXC+lhcA29ZBXYD9hOMbmFz7tE16TKLcMrRNWhDWKbwOVIZjyM
A6Wywtr1XudycnsbEZT8XPkVR67AC627U7uGnEsreLp6TfS315ehSbBAm2/c0fZBSYPwN7UQ4x5x
gAac9EuyXYf/K9bLsBKgAo4uDNAPSK6ndrdTygsgF1zpTzTWxY1GlCG3oUJIp9YME+wAS+9Du+CX
gc4Bvc20eZYrkisQfJjSysA+yA7voea6ulpLe8haC2CRQX9KJdrfeXW2tZlRd+RNTouxwqyIlQlE
RgE8ge/duBOWkzj2njjaXiHqY7dOFcdG16hxgq9SFxE6meE3P6z68MV/HtZT4vJbO9naJU7OpNyT
szsiZz1rAYDuHjIVCQwmwxxgkrMvIOf6IXb1njZDKf+EUiHkMFsDgoEj9RsIBPK8ifCLRrNdTSoe
3HTj9fFTBLwRlXFtUI/l3LRQyn8HchyinVzk8NQsY8XKBw==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity watch_events_int is
port(
  Data :  in std_logic_vector(71 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(71 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end watch_events_int;
architecture beh of watch_events_int is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo_sc.watch_events_int\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(71 downto 0);
  Full: out std_logic;
  Empty: out std_logic;
  Q : out std_logic_vector(71 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_inst: \~fifo_sc.watch_events_int\
port map(
  Clk => Clk,
  Reset => Reset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(71 downto 0) => Data(71 downto 0),
  Full => NN_0,
  Empty => NN,
  Q(71 downto 0) => Q(71 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
